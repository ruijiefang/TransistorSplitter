.SUBCKT DFFLQNx3_ASAP7_75t_L CLK D QN VDD VSS
MM27 clkb clkn VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MM0 clkn CLK VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MM24 QN SH VSS VSS nmos_lvt w=243.00n l=20n nfin=9
MM17 SH clkb pd5 VSS nmos_lvt w=27.0n l=20n nfin=1
MM16 pd5 SS VSS VSS nmos_lvt w=27.0n l=20n nfin=1
MM14 SS SH VSS VSS nmos_lvt w=27.0n l=20n nfin=1
MM12 MS clkn SH VSS nmos_lvt w=27.0n l=20n nfin=1
MM6 MS MH VSS VSS nmos_lvt w=27.0n l=20n nfin=1
MM9 MH clkn pd3 VSS nmos_lvt w=27.0n l=20n nfin=1
MM8 pd3 MS VSS VSS nmos_lvt w=27.0n l=20n nfin=1
MM5 pd1 D VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM4 MH clkb pd1 VSS nmos_lvt w=81.0n l=20n nfin=3
MM26 clkb clkn VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MM2 clkn CLK VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MM25 QN SH VDD VDD pmos_lvt w=243.00n l=20n nfin=9
MM19 pd4 SS VDD VDD pmos_lvt w=27n l=20n nfin=1
MM18 SH clkn pd4 VDD pmos_lvt w=27n l=20n nfin=1
MM15 SS SH VDD VDD pmos_lvt w=27n l=20n nfin=1
MM13 MS clkb SH VDD pmos_lvt w=27n l=20n nfin=1
MM7 MS MH VDD VDD pmos_lvt w=27n l=20n nfin=1
MM11 pd2 MS VDD VDD pmos_lvt w=27n l=20n nfin=1
MM10 MH clkb pd2 VDD pmos_lvt w=27n l=20n nfin=1
MM1 MH clkn pu1 VDD pmos_lvt w=81.0n l=20n nfin=3
MM3 pu1 D VDD VDD pmos_lvt w=81.0n l=20n nfin=3
.ENDS

