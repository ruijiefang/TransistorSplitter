.SUBCKT DLLx3_ASAP7_75t_L CLK D Q VDD VSS
MM24 Q MH VSS VSS nmos_lvt w=243.00n l=20n nfin=9
MM6 net30 MH VSS VSS nmos_lvt w=27.0n l=20n nfin=1
MM9 MH clkb pd3 VSS nmos_lvt w=27.0n l=20n nfin=1
MM8 pd3 net30 VSS VSS nmos_lvt w=27.0n l=20n nfin=1
MM23 clkb clkn VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MM5 pd1 D VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM4 MH clkn pd1 VSS nmos_lvt w=81.0n l=20n nfin=3
MM20 clkn CLK VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MM25 Q MH VDD VDD pmos_lvt w=243.00n l=20n nfin=9
MM7 net30 MH VDD VDD pmos_lvt w=27n l=20n nfin=1
MM11 pd2 net30 VDD VDD pmos_lvt w=27n l=20n nfin=1
MM10 MH clkn pd2 VDD pmos_lvt w=27n l=20n nfin=1
MM22 clkb clkn VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MM1 MH clkb pu1 VDD pmos_lvt w=81.0n l=20n nfin=3
MM3 pu1 D VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM21 clkn CLK VDD VDD pmos_lvt w=54.0n l=20n nfin=2
.ENDS
