.SUBCKT FAx1_ASAP7_75t_L A B CI CON SN VDD VSS
MM22 SN CI net081 VDD pmos_lvt w=81.0n l=20n nfin=3
MM21 net081 B net082 VDD pmos_lvt w=81.0n l=20n nfin=3
MM20 net082 A VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM15 SN CON net027 VDD pmos_lvt w=81.0n l=20n nfin=3
MM14 net027 CI VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM13 net027 B VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM12 net027 A VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM5 CON A net37 VDD pmos_lvt w=81.0n l=20n nfin=3
MM6 net37 B VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM2 net27 B VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM1 CON CI net27 VDD pmos_lvt w=81.0n l=20n nfin=3
MM0 net27 A VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM25 SN CI net080 VSS nmos_lvt w=81.0n l=20n nfin=3
MM24 net080 B net079 VSS nmos_lvt w=81.0n l=20n nfin=3
MM23 net079 A VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM19 VSS CI net067 VSS nmos_lvt w=81.0n l=20n nfin=3
MM18 VSS B net067 VSS nmos_lvt w=81.0n l=20n nfin=3
MM17 VSS A net067 VSS nmos_lvt w=81.0n l=20n nfin=3
MM16 net067 CON SN VSS nmos_lvt w=81.0n l=20n nfin=3
MM11 VSS B net25 VSS nmos_lvt w=81.0n l=20n nfin=3
MM10 VSS B net36 VSS nmos_lvt w=81.0n l=20n nfin=3
MM9 VSS A net25 VSS nmos_lvt w=81.0n l=20n nfin=3
MM8 net36 A CON VSS nmos_lvt w=81.0n l=20n nfin=3
MM7 net25 CI CON VSS nmos_lvt w=81.0n l=20n nfin=3
.ENDS

