.SUBCKT adder8 a_7_ a_6_ a_5_ a_4_ a_3_ a_2_ a_1_ a_0_ b_7_ b_6_ b_5_ b_4_ b_3_ b_2_ b_1_ b_0_ y_7_ y_6_ y_5_ y_4_ y_3_ y_2_ y_1_ y_0_
* FAxp33_ASAP7_6t_L add_4_U1_0
MMP0_add_4_U1_0_inst0_MM22 n18 add_4_CI inst0_net081 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP1_add_4_U1_0_inst0_MM21 inst0_net081 b_0_ inst0_net082 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP2_add_4_U1_0_inst0_MM20 inst0_net082 a_0_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP3_add_4_U1_0_inst0_MM15 n18 n19 inst0_net027 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP4_add_4_U1_0_inst0_MM14 inst0_net027 add_4_CI VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP5_add_4_U1_0_inst0_MM13 inst0_net027 b_0_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP6_add_4_U1_0_inst0_MM12 inst0_net027 a_0_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP7_add_4_U1_0_inst0_MM5 n19 a_0_ inst0_net37 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP8_add_4_U1_0_inst0_MM6 inst0_net37 b_0_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP9_add_4_U1_0_inst0_MM2 inst0_net27 b_0_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP10_add_4_U1_0_inst0_MM1 n19 add_4_CI inst0_net27 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP11_add_4_U1_0_inst0_MM0 inst0_net27 a_0_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMN12_add_4_U1_0_inst0_MM25 n18 add_4_CI inst0_net080 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN13_add_4_U1_0_inst0_MM24 inst0_net080 b_0_ inst0_net079 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN14_add_4_U1_0_inst0_MM23 inst0_net079 a_0_ VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MMN15_add_4_U1_0_inst0_MM19 VSS add_4_CI inst0_net067 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN16_add_4_U1_0_inst0_MM18 VSS b_0_ inst0_net067 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN17_add_4_U1_0_inst0_MM17 VSS a_0_ inst0_net067 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN18_add_4_U1_0_inst0_MM16 inst0_net067 n19 n18 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN19_add_4_U1_0_inst0_MM11 VSS b_0_ inst0_net25 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN20_add_4_U1_0_inst0_MM10 VSS b_0_ inst0_net36 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN21_add_4_U1_0_inst0_MM9 VSS a_0_ inst0_net25 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN22_add_4_U1_0_inst0_MM8 inst0_net36 a_0_ n19 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN23_add_4_U1_0_inst0_MM7 inst0_net25 add_4_CI n19 VSS nmos_lvt w=54.0n l=20n nfin=2
* FAxp33_ASAP7_6t_L add_4_U1_1
MMP24_add_4_U1_1_inst1_MM22 n20 n16 inst1_net081 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP25_add_4_U1_1_inst1_MM21 inst1_net081 b_1_ inst1_net082 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP26_add_4_U1_1_inst1_MM20 inst1_net082 a_1_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP27_add_4_U1_1_inst1_MM15 n20 n21 inst1_net027 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP28_add_4_U1_1_inst1_MM14 inst1_net027 n16 VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP29_add_4_U1_1_inst1_MM13 inst1_net027 b_1_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP30_add_4_U1_1_inst1_MM12 inst1_net027 a_1_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP31_add_4_U1_1_inst1_MM5 n21 a_1_ inst1_net37 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP32_add_4_U1_1_inst1_MM6 inst1_net37 b_1_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP33_add_4_U1_1_inst1_MM2 inst1_net27 b_1_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP34_add_4_U1_1_inst1_MM1 n21 n16 inst1_net27 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP35_add_4_U1_1_inst1_MM0 inst1_net27 a_1_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMN36_add_4_U1_1_inst1_MM25 n20 n16 inst1_net080 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN37_add_4_U1_1_inst1_MM24 inst1_net080 b_1_ inst1_net079 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN38_add_4_U1_1_inst1_MM23 inst1_net079 a_1_ VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MMN39_add_4_U1_1_inst1_MM19 VSS n16 inst1_net067 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN40_add_4_U1_1_inst1_MM18 VSS b_1_ inst1_net067 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN41_add_4_U1_1_inst1_MM17 VSS a_1_ inst1_net067 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN42_add_4_U1_1_inst1_MM16 inst1_net067 n21 n20 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN43_add_4_U1_1_inst1_MM11 VSS b_1_ inst1_net25 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN44_add_4_U1_1_inst1_MM10 VSS b_1_ inst1_net36 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN45_add_4_U1_1_inst1_MM9 VSS a_1_ inst1_net25 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN46_add_4_U1_1_inst1_MM8 inst1_net36 a_1_ n21 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN47_add_4_U1_1_inst1_MM7 inst1_net25 n16 n21 VSS nmos_lvt w=54.0n l=20n nfin=2
* FAxp33_ASAP7_6t_L add_4_U1_2
MMP48_add_4_U1_2_inst2_MM22 n22 n14 inst2_net081 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP49_add_4_U1_2_inst2_MM21 inst2_net081 b_2_ inst2_net082 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP50_add_4_U1_2_inst2_MM20 inst2_net082 a_2_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP51_add_4_U1_2_inst2_MM15 n22 n23 inst2_net027 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP52_add_4_U1_2_inst2_MM14 inst2_net027 n14 VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP53_add_4_U1_2_inst2_MM13 inst2_net027 b_2_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP54_add_4_U1_2_inst2_MM12 inst2_net027 a_2_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP55_add_4_U1_2_inst2_MM5 n23 a_2_ inst2_net37 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP56_add_4_U1_2_inst2_MM6 inst2_net37 b_2_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP57_add_4_U1_2_inst2_MM2 inst2_net27 b_2_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP58_add_4_U1_2_inst2_MM1 n23 n14 inst2_net27 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP59_add_4_U1_2_inst2_MM0 inst2_net27 a_2_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMN60_add_4_U1_2_inst2_MM25 n22 n14 inst2_net080 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN61_add_4_U1_2_inst2_MM24 inst2_net080 b_2_ inst2_net079 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN62_add_4_U1_2_inst2_MM23 inst2_net079 a_2_ VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MMN63_add_4_U1_2_inst2_MM19 VSS n14 inst2_net067 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN64_add_4_U1_2_inst2_MM18 VSS b_2_ inst2_net067 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN65_add_4_U1_2_inst2_MM17 VSS a_2_ inst2_net067 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN66_add_4_U1_2_inst2_MM16 inst2_net067 n23 n22 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN67_add_4_U1_2_inst2_MM11 VSS b_2_ inst2_net25 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN68_add_4_U1_2_inst2_MM10 VSS b_2_ inst2_net36 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN69_add_4_U1_2_inst2_MM9 VSS a_2_ inst2_net25 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN70_add_4_U1_2_inst2_MM8 inst2_net36 a_2_ n23 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN71_add_4_U1_2_inst2_MM7 inst2_net25 n14 n23 VSS nmos_lvt w=54.0n l=20n nfin=2
* FAxp33_ASAP7_6t_L add_4_U1_3
MMP72_add_4_U1_3_inst3_MM22 n24 n12 inst3_net081 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP73_add_4_U1_3_inst3_MM21 inst3_net081 b_3_ inst3_net082 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP74_add_4_U1_3_inst3_MM20 inst3_net082 a_3_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP75_add_4_U1_3_inst3_MM15 n24 n25 inst3_net027 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP76_add_4_U1_3_inst3_MM14 inst3_net027 n12 VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP77_add_4_U1_3_inst3_MM13 inst3_net027 b_3_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP78_add_4_U1_3_inst3_MM12 inst3_net027 a_3_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP79_add_4_U1_3_inst3_MM5 n25 a_3_ inst3_net37 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP80_add_4_U1_3_inst3_MM6 inst3_net37 b_3_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP81_add_4_U1_3_inst3_MM2 inst3_net27 b_3_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP82_add_4_U1_3_inst3_MM1 n25 n12 inst3_net27 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP83_add_4_U1_3_inst3_MM0 inst3_net27 a_3_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMN84_add_4_U1_3_inst3_MM25 n24 n12 inst3_net080 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN85_add_4_U1_3_inst3_MM24 inst3_net080 b_3_ inst3_net079 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN86_add_4_U1_3_inst3_MM23 inst3_net079 a_3_ VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MMN87_add_4_U1_3_inst3_MM19 VSS n12 inst3_net067 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN88_add_4_U1_3_inst3_MM18 VSS b_3_ inst3_net067 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN89_add_4_U1_3_inst3_MM17 VSS a_3_ inst3_net067 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN90_add_4_U1_3_inst3_MM16 inst3_net067 n25 n24 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN91_add_4_U1_3_inst3_MM11 VSS b_3_ inst3_net25 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN92_add_4_U1_3_inst3_MM10 VSS b_3_ inst3_net36 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN93_add_4_U1_3_inst3_MM9 VSS a_3_ inst3_net25 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN94_add_4_U1_3_inst3_MM8 inst3_net36 a_3_ n25 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN95_add_4_U1_3_inst3_MM7 inst3_net25 n12 n25 VSS nmos_lvt w=54.0n l=20n nfin=2
* FAxp33_ASAP7_6t_L add_4_U1_4
MMP96_add_4_U1_4_inst4_MM22 n26 n10 inst4_net081 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP97_add_4_U1_4_inst4_MM21 inst4_net081 b_4_ inst4_net082 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP98_add_4_U1_4_inst4_MM20 inst4_net082 a_4_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP99_add_4_U1_4_inst4_MM15 n26 n27 inst4_net027 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP100_add_4_U1_4_inst4_MM14 inst4_net027 n10 VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP101_add_4_U1_4_inst4_MM13 inst4_net027 b_4_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP102_add_4_U1_4_inst4_MM12 inst4_net027 a_4_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP103_add_4_U1_4_inst4_MM5 n27 a_4_ inst4_net37 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP104_add_4_U1_4_inst4_MM6 inst4_net37 b_4_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP105_add_4_U1_4_inst4_MM2 inst4_net27 b_4_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP106_add_4_U1_4_inst4_MM1 n27 n10 inst4_net27 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP107_add_4_U1_4_inst4_MM0 inst4_net27 a_4_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMN108_add_4_U1_4_inst4_MM25 n26 n10 inst4_net080 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN109_add_4_U1_4_inst4_MM24 inst4_net080 b_4_ inst4_net079 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN110_add_4_U1_4_inst4_MM23 inst4_net079 a_4_ VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MMN111_add_4_U1_4_inst4_MM19 VSS n10 inst4_net067 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN112_add_4_U1_4_inst4_MM18 VSS b_4_ inst4_net067 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN113_add_4_U1_4_inst4_MM17 VSS a_4_ inst4_net067 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN114_add_4_U1_4_inst4_MM16 inst4_net067 n27 n26 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN115_add_4_U1_4_inst4_MM11 VSS b_4_ inst4_net25 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN116_add_4_U1_4_inst4_MM10 VSS b_4_ inst4_net36 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN117_add_4_U1_4_inst4_MM9 VSS a_4_ inst4_net25 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN118_add_4_U1_4_inst4_MM8 inst4_net36 a_4_ n27 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN119_add_4_U1_4_inst4_MM7 inst4_net25 n10 n27 VSS nmos_lvt w=54.0n l=20n nfin=2
* FAxp33_ASAP7_6t_L add_4_U1_5
MMP120_add_4_U1_5_inst5_MM22 n28 n8 inst5_net081 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP121_add_4_U1_5_inst5_MM21 inst5_net081 b_5_ inst5_net082 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP122_add_4_U1_5_inst5_MM20 inst5_net082 a_5_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP123_add_4_U1_5_inst5_MM15 n28 n29 inst5_net027 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP124_add_4_U1_5_inst5_MM14 inst5_net027 n8 VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP125_add_4_U1_5_inst5_MM13 inst5_net027 b_5_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP126_add_4_U1_5_inst5_MM12 inst5_net027 a_5_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP127_add_4_U1_5_inst5_MM5 n29 a_5_ inst5_net37 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP128_add_4_U1_5_inst5_MM6 inst5_net37 b_5_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP129_add_4_U1_5_inst5_MM2 inst5_net27 b_5_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP130_add_4_U1_5_inst5_MM1 n29 n8 inst5_net27 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP131_add_4_U1_5_inst5_MM0 inst5_net27 a_5_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMN132_add_4_U1_5_inst5_MM25 n28 n8 inst5_net080 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN133_add_4_U1_5_inst5_MM24 inst5_net080 b_5_ inst5_net079 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN134_add_4_U1_5_inst5_MM23 inst5_net079 a_5_ VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MMN135_add_4_U1_5_inst5_MM19 VSS n8 inst5_net067 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN136_add_4_U1_5_inst5_MM18 VSS b_5_ inst5_net067 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN137_add_4_U1_5_inst5_MM17 VSS a_5_ inst5_net067 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN138_add_4_U1_5_inst5_MM16 inst5_net067 n29 n28 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN139_add_4_U1_5_inst5_MM11 VSS b_5_ inst5_net25 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN140_add_4_U1_5_inst5_MM10 VSS b_5_ inst5_net36 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN141_add_4_U1_5_inst5_MM9 VSS a_5_ inst5_net25 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN142_add_4_U1_5_inst5_MM8 inst5_net36 a_5_ n29 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN143_add_4_U1_5_inst5_MM7 inst5_net25 n8 n29 VSS nmos_lvt w=54.0n l=20n nfin=2
* FAxp33_ASAP7_6t_L add_4_U1_6
MMP144_add_4_U1_6_inst6_MM22 n30 n6 inst6_net081 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP145_add_4_U1_6_inst6_MM21 inst6_net081 b_6_ inst6_net082 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP146_add_4_U1_6_inst6_MM20 inst6_net082 a_6_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP147_add_4_U1_6_inst6_MM15 n30 n31 inst6_net027 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP148_add_4_U1_6_inst6_MM14 inst6_net027 n6 VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP149_add_4_U1_6_inst6_MM13 inst6_net027 b_6_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP150_add_4_U1_6_inst6_MM12 inst6_net027 a_6_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP151_add_4_U1_6_inst6_MM5 n31 a_6_ inst6_net37 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP152_add_4_U1_6_inst6_MM6 inst6_net37 b_6_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP153_add_4_U1_6_inst6_MM2 inst6_net27 b_6_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP154_add_4_U1_6_inst6_MM1 n31 n6 inst6_net27 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP155_add_4_U1_6_inst6_MM0 inst6_net27 a_6_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMN156_add_4_U1_6_inst6_MM25 n30 n6 inst6_net080 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN157_add_4_U1_6_inst6_MM24 inst6_net080 b_6_ inst6_net079 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN158_add_4_U1_6_inst6_MM23 inst6_net079 a_6_ VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MMN159_add_4_U1_6_inst6_MM19 VSS n6 inst6_net067 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN160_add_4_U1_6_inst6_MM18 VSS b_6_ inst6_net067 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN161_add_4_U1_6_inst6_MM17 VSS a_6_ inst6_net067 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN162_add_4_U1_6_inst6_MM16 inst6_net067 n31 n30 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN163_add_4_U1_6_inst6_MM11 VSS b_6_ inst6_net25 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN164_add_4_U1_6_inst6_MM10 VSS b_6_ inst6_net36 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN165_add_4_U1_6_inst6_MM9 VSS a_6_ inst6_net25 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN166_add_4_U1_6_inst6_MM8 inst6_net36 a_6_ n31 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN167_add_4_U1_6_inst6_MM7 inst6_net25 n6 n31 VSS nmos_lvt w=54.0n l=20n nfin=2

* FAxp33_ASAP7_6t_L add_4_U1_7
MMP168_add_4_U1_7_inst7_MM22 n32 n4 inst7_net081 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP169_add_4_U1_7_inst7_MM21 inst7_net081 b_7_ inst7_net082 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP170_add_4_U1_7_inst7_MM20 inst7_net082 a_7_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP171_add_4_U1_7_inst7_MM15 n32 inst7_CON inst7_net027 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP172_add_4_U1_7_inst7_MM14 inst7_net027 n4 VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP173_add_4_U1_7_inst7_MM13 inst7_net027 b_7_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP174_add_4_U1_7_inst7_MM12 inst7_net027 a_7_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP175_add_4_U1_7_inst7_MM5 inst7_CON a_7_ inst7_net37 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP176_add_4_U1_7_inst7_MM6 inst7_net37 b_7_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP177_add_4_U1_7_inst7_MM2 inst7_net27 b_7_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP178_add_4_U1_7_inst7_MM1 inst7_CON n4 inst7_net27 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP179_add_4_U1_7_inst7_MM0 inst7_net27 a_7_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMN180_add_4_U1_7_inst7_MM25 n32 n4 inst7_net080 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN181_add_4_U1_7_inst7_MM24 inst7_net080 b_7_ inst7_net079 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN182_add_4_U1_7_inst7_MM23 inst7_net079 a_7_ VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MMN183_add_4_U1_7_inst7_MM19 VSS n4 inst7_net067 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN184_add_4_U1_7_inst7_MM18 VSS b_7_ inst7_net067 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN185_add_4_U1_7_inst7_MM17 VSS a_7_ inst7_net067 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN186_add_4_U1_7_inst7_MM16 inst7_net067 inst7_CON n32 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN187_add_4_U1_7_inst7_MM11 VSS b_7_ inst7_net25 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN188_add_4_U1_7_inst7_MM10 VSS b_7_ inst7_net36 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN189_add_4_U1_7_inst7_MM9 VSS a_7_ inst7_net25 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN190_add_4_U1_7_inst7_MM8 inst7_net36 a_7_ inst7_CON VSS nmos_lvt w=54.0n l=20n nfin=2
MMN191_add_4_U1_7_inst7_MM7 inst7_net25 n4 inst7_CON VSS nmos_lvt w=54.0n l=20n nfin=2
* TIELOxp5_ASAP7_6t_L U3
MMP192_U3_inst8_MM1 inst8_net9 add_4_CI VDD VDD pmos_lvt w=27.0n l=20n nfin=1
MMN193_U3_inst8_MM2 add_4_CI inst8_net9 VSS VSS nmos_lvt w=27.0n l=20n nfin=1
* INVx1_ASAP7_6t_L U4
MMN194_U4_inst9_MM0 y_7_ n32 VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MMP195_U4_inst9_MM1 y_7_ n32 VDD VDD pmos_lvt w=54.0n l=20n nfin=2
* INVx1_ASAP7_6t_L U5
MMN196_U5_inst10_MM0 n4 n31 VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MMP197_U5_inst10_MM1 n4 n31 VDD VDD pmos_lvt w=54.0n l=20n nfin=2
* INVx1_ASAP7_6t_L U6
MMN198_U6_inst11_MM0 y_6_ n30 VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MMP199_U6_inst11_MM1 y_6_ n30 VDD VDD pmos_lvt w=54.0n l=20n nfin=2
* INVx1_ASAP7_6t_L U7
MMN200_U7_inst12_MM0 n6 n29 VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MMP201_U7_inst12_MM1 n6 n29 VDD VDD pmos_lvt w=54.0n l=20n nfin=2
* INVx1_ASAP7_6t_L U8
MMN202_U8_inst13_MM0 y_5_ n28 VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MMP203_U8_inst13_MM1 y_5_ n28 VDD VDD pmos_lvt w=54.0n l=20n nfin=2
* INVx1_ASAP7_6t_L U9
MMN204_U9_inst14_MM0 n8 n27 VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MMP205_U9_inst14_MM1 n8 n27 VDD VDD pmos_lvt w=54.0n l=20n nfin=2
* INVx1_ASAP7_6t_L U10
MMN206_U10_inst15_MM0 y_4_ n26 VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MMP207_U10_inst15_MM1 y_4_ n26 VDD VDD pmos_lvt w=54.0n l=20n nfin=2
* INVx1_ASAP7_6t_L U11
MMN208_U11_inst16_MM0 n10 n25 VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MMP209_U11_inst16_MM1 n10 n25 VDD VDD pmos_lvt w=54.0n l=20n nfin=2
* INVx1_ASAP7_6t_L U12
MMN210_U12_inst17_MM0 y_3_ n24 VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MMP211_U12_inst17_MM1 y_3_ n24 VDD VDD pmos_lvt w=54.0n l=20n nfin=2
* INVx1_ASAP7_6t_L U13
MMN212_U13_inst18_MM0 n12 n23 VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MMP213_U13_inst18_MM1 n12 n23 VDD VDD pmos_lvt w=54.0n l=20n nfin=2
* INVx1_ASAP7_6t_L U14
MMN214_U14_inst19_MM0 y_2_ n22 VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MMP215_U14_inst19_MM1 y_2_ n22 VDD VDD pmos_lvt w=54.0n l=20n nfin=2
* INVx1_ASAP7_6t_L U15
MMN216_U15_inst20_MM0 n14 n21 VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MMP217_U15_inst20_MM1 n14 n21 VDD VDD pmos_lvt w=54.0n l=20n nfin=2
* INVx1_ASAP7_6t_L U16
MMN218_U16_inst21_MM0 y_1_ n20 VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MMP219_U16_inst21_MM1 y_1_ n20 VDD VDD pmos_lvt w=54.0n l=20n nfin=2
* INVx1_ASAP7_6t_L U17
MMN220_U17_inst22_MM0 n16 n19 VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MMP221_U17_inst22_MM1 n16 n19 VDD VDD pmos_lvt w=54.0n l=20n nfin=2
* INVx1_ASAP7_6t_L U18
MMN222_U18_inst23_MM0 y_0_ n18 VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MMP223_U18_inst23_MM1 y_0_ n18 VDD VDD pmos_lvt w=54.0n l=20n nfin=2
.ENDS
