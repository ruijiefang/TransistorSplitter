.SUBCKT mul4x4 a_3_ a_2_ a_1_ a_0_ b_3_ b_2_ b_1_ b_0_ y_7_ y_6_ y_5_ y_4_ y_3_ y_2_ y_1_ y_0_


* FAxp33_ASAP7_6t_L dp_cluster_0_mult_4_S3_2_2
MMP0_dp_cluster_0_mult_4_S3_2_2_inst0_MM22 n39 dp_cluster_0_mult_4_ab_1__3_ inst0_net081 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP1_dp_cluster_0_mult_4_S3_2_2_inst0_MM21 inst0_net081 n7 inst0_net082 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP2_dp_cluster_0_mult_4_S3_2_2_inst0_MM20 inst0_net082 dp_cluster_0_mult_4_ab_2__2_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP3_dp_cluster_0_mult_4_S3_2_2_inst0_MM15 n39 n40 inst0_net027 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP4_dp_cluster_0_mult_4_S3_2_2_inst0_MM14 inst0_net027 dp_cluster_0_mult_4_ab_1__3_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP5_dp_cluster_0_mult_4_S3_2_2_inst0_MM13 inst0_net027 n7 VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP6_dp_cluster_0_mult_4_S3_2_2_inst0_MM12 inst0_net027 dp_cluster_0_mult_4_ab_2__2_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP7_dp_cluster_0_mult_4_S3_2_2_inst0_MM5 n40 dp_cluster_0_mult_4_ab_2__2_ inst0_net37 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP8_dp_cluster_0_mult_4_S3_2_2_inst0_MM6 inst0_net37 n7 VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP9_dp_cluster_0_mult_4_S3_2_2_inst0_MM2 inst0_net27 n7 VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP10_dp_cluster_0_mult_4_S3_2_2_inst0_MM1 n40 dp_cluster_0_mult_4_ab_1__3_ inst0_net27 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP11_dp_cluster_0_mult_4_S3_2_2_inst0_MM0 inst0_net27 dp_cluster_0_mult_4_ab_2__2_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMN12_dp_cluster_0_mult_4_S3_2_2_inst0_MM25 n39 dp_cluster_0_mult_4_ab_1__3_ inst0_net080 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN13_dp_cluster_0_mult_4_S3_2_2_inst0_MM24 inst0_net080 n7 inst0_net079 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN14_dp_cluster_0_mult_4_S3_2_2_inst0_MM23 inst0_net079 dp_cluster_0_mult_4_ab_2__2_ VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MMN15_dp_cluster_0_mult_4_S3_2_2_inst0_MM19 VSS dp_cluster_0_mult_4_ab_1__3_ inst0_net067 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN16_dp_cluster_0_mult_4_S3_2_2_inst0_MM18 VSS n7 inst0_net067 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN17_dp_cluster_0_mult_4_S3_2_2_inst0_MM17 VSS dp_cluster_0_mult_4_ab_2__2_ inst0_net067 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN18_dp_cluster_0_mult_4_S3_2_2_inst0_MM16 inst0_net067 n40 n39 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN19_dp_cluster_0_mult_4_S3_2_2_inst0_MM11 VSS n7 inst0_net25 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN20_dp_cluster_0_mult_4_S3_2_2_inst0_MM10 VSS n7 inst0_net36 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN21_dp_cluster_0_mult_4_S3_2_2_inst0_MM9 VSS dp_cluster_0_mult_4_ab_2__2_ inst0_net25 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN22_dp_cluster_0_mult_4_S3_2_2_inst0_MM8 inst0_net36 dp_cluster_0_mult_4_ab_2__2_ n40 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN23_dp_cluster_0_mult_4_S3_2_2_inst0_MM7 inst0_net25 dp_cluster_0_mult_4_ab_1__3_ n40 VSS nmos_lvt w=54.0n l=20n nfin=2

* FAxp33_ASAP7_6t_L dp_cluster_0_mult_4_S2_2_1
MMP24_dp_cluster_0_mult_4_S2_2_1_inst1_MM22 n41 n9 inst1_net081 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP25_dp_cluster_0_mult_4_S2_2_1_inst1_MM21 inst1_net081 n4 inst1_net082 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP26_dp_cluster_0_mult_4_S2_2_1_inst1_MM20 inst1_net082 dp_cluster_0_mult_4_ab_2__1_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP27_dp_cluster_0_mult_4_S2_2_1_inst1_MM15 n41 n42 inst1_net027 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP28_dp_cluster_0_mult_4_S2_2_1_inst1_MM14 inst1_net027 n9 VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP29_dp_cluster_0_mult_4_S2_2_1_inst1_MM13 inst1_net027 n4 VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP30_dp_cluster_0_mult_4_S2_2_1_inst1_MM12 inst1_net027 dp_cluster_0_mult_4_ab_2__1_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP31_dp_cluster_0_mult_4_S2_2_1_inst1_MM5 n42 dp_cluster_0_mult_4_ab_2__1_ inst1_net37 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP32_dp_cluster_0_mult_4_S2_2_1_inst1_MM6 inst1_net37 n4 VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP33_dp_cluster_0_mult_4_S2_2_1_inst1_MM2 inst1_net27 n4 VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP34_dp_cluster_0_mult_4_S2_2_1_inst1_MM1 n42 n9 inst1_net27 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP35_dp_cluster_0_mult_4_S2_2_1_inst1_MM0 inst1_net27 dp_cluster_0_mult_4_ab_2__1_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMN36_dp_cluster_0_mult_4_S2_2_1_inst1_MM25 n41 n9 inst1_net080 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN37_dp_cluster_0_mult_4_S2_2_1_inst1_MM24 inst1_net080 n4 inst1_net079 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN38_dp_cluster_0_mult_4_S2_2_1_inst1_MM23 inst1_net079 dp_cluster_0_mult_4_ab_2__1_ VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MMN39_dp_cluster_0_mult_4_S2_2_1_inst1_MM19 VSS n9 inst1_net067 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN40_dp_cluster_0_mult_4_S2_2_1_inst1_MM18 VSS n4 inst1_net067 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN41_dp_cluster_0_mult_4_S2_2_1_inst1_MM17 VSS dp_cluster_0_mult_4_ab_2__1_ inst1_net067 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN42_dp_cluster_0_mult_4_S2_2_1_inst1_MM16 inst1_net067 n42 n41 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN43_dp_cluster_0_mult_4_S2_2_1_inst1_MM11 VSS n4 inst1_net25 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN44_dp_cluster_0_mult_4_S2_2_1_inst1_MM10 VSS n4 inst1_net36 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN45_dp_cluster_0_mult_4_S2_2_1_inst1_MM9 VSS dp_cluster_0_mult_4_ab_2__1_ inst1_net25 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN46_dp_cluster_0_mult_4_S2_2_1_inst1_MM8 inst1_net36 dp_cluster_0_mult_4_ab_2__1_ n42 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN47_dp_cluster_0_mult_4_S2_2_1_inst1_MM7 inst1_net25 n9 n42 VSS nmos_lvt w=54.0n l=20n nfin=2

* FAxp33_ASAP7_6t_L dp_cluster_0_mult_4_S1_2_0
MMP48_dp_cluster_0_mult_4_S1_2_0_inst2_MM22 n43 n8 inst2_net081 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP49_dp_cluster_0_mult_4_S1_2_0_inst2_MM21 inst2_net081 n3 inst2_net082 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP50_dp_cluster_0_mult_4_S1_2_0_inst2_MM20 inst2_net082 dp_cluster_0_mult_4_ab_2__0_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP51_dp_cluster_0_mult_4_S1_2_0_inst2_MM15 n43 n44 inst2_net027 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP52_dp_cluster_0_mult_4_S1_2_0_inst2_MM14 inst2_net027 n8 VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP53_dp_cluster_0_mult_4_S1_2_0_inst2_MM13 inst2_net027 n3 VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP54_dp_cluster_0_mult_4_S1_2_0_inst2_MM12 inst2_net027 dp_cluster_0_mult_4_ab_2__0_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP55_dp_cluster_0_mult_4_S1_2_0_inst2_MM5 n44 dp_cluster_0_mult_4_ab_2__0_ inst2_net37 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP56_dp_cluster_0_mult_4_S1_2_0_inst2_MM6 inst2_net37 n3 VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP57_dp_cluster_0_mult_4_S1_2_0_inst2_MM2 inst2_net27 n3 VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP58_dp_cluster_0_mult_4_S1_2_0_inst2_MM1 n44 n8 inst2_net27 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP59_dp_cluster_0_mult_4_S1_2_0_inst2_MM0 inst2_net27 dp_cluster_0_mult_4_ab_2__0_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMN60_dp_cluster_0_mult_4_S1_2_0_inst2_MM25 n43 n8 inst2_net080 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN61_dp_cluster_0_mult_4_S1_2_0_inst2_MM24 inst2_net080 n3 inst2_net079 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN62_dp_cluster_0_mult_4_S1_2_0_inst2_MM23 inst2_net079 dp_cluster_0_mult_4_ab_2__0_ VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MMN63_dp_cluster_0_mult_4_S1_2_0_inst2_MM19 VSS n8 inst2_net067 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN64_dp_cluster_0_mult_4_S1_2_0_inst2_MM18 VSS n3 inst2_net067 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN65_dp_cluster_0_mult_4_S1_2_0_inst2_MM17 VSS dp_cluster_0_mult_4_ab_2__0_ inst2_net067 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN66_dp_cluster_0_mult_4_S1_2_0_inst2_MM16 inst2_net067 n44 n43 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN67_dp_cluster_0_mult_4_S1_2_0_inst2_MM11 VSS n3 inst2_net25 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN68_dp_cluster_0_mult_4_S1_2_0_inst2_MM10 VSS n3 inst2_net36 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN69_dp_cluster_0_mult_4_S1_2_0_inst2_MM9 VSS dp_cluster_0_mult_4_ab_2__0_ inst2_net25 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN70_dp_cluster_0_mult_4_S1_2_0_inst2_MM8 inst2_net36 dp_cluster_0_mult_4_ab_2__0_ n44 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN71_dp_cluster_0_mult_4_S1_2_0_inst2_MM7 inst2_net25 n8 n44 VSS nmos_lvt w=54.0n l=20n nfin=2

* FAxp33_ASAP7_6t_L dp_cluster_0_mult_4_S5_2
MMP72_dp_cluster_0_mult_4_S5_2_inst3_MM22 n45 dp_cluster_0_mult_4_ab_2__3_ inst3_net081 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP73_dp_cluster_0_mult_4_S5_2_inst3_MM21 inst3_net081 n30 inst3_net082 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP74_dp_cluster_0_mult_4_S5_2_inst3_MM20 inst3_net082 dp_cluster_0_mult_4_ab_3__2_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP75_dp_cluster_0_mult_4_S5_2_inst3_MM15 n45 n46 inst3_net027 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP76_dp_cluster_0_mult_4_S5_2_inst3_MM14 inst3_net027 dp_cluster_0_mult_4_ab_2__3_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP77_dp_cluster_0_mult_4_S5_2_inst3_MM13 inst3_net027 n30 VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP78_dp_cluster_0_mult_4_S5_2_inst3_MM12 inst3_net027 dp_cluster_0_mult_4_ab_3__2_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP79_dp_cluster_0_mult_4_S5_2_inst3_MM5 n46 dp_cluster_0_mult_4_ab_3__2_ inst3_net37 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP80_dp_cluster_0_mult_4_S5_2_inst3_MM6 inst3_net37 n30 VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP81_dp_cluster_0_mult_4_S5_2_inst3_MM2 inst3_net27 n30 VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP82_dp_cluster_0_mult_4_S5_2_inst3_MM1 n46 dp_cluster_0_mult_4_ab_2__3_ inst3_net27 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP83_dp_cluster_0_mult_4_S5_2_inst3_MM0 inst3_net27 dp_cluster_0_mult_4_ab_3__2_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMN84_dp_cluster_0_mult_4_S5_2_inst3_MM25 n45 dp_cluster_0_mult_4_ab_2__3_ inst3_net080 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN85_dp_cluster_0_mult_4_S5_2_inst3_MM24 inst3_net080 n30 inst3_net079 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN86_dp_cluster_0_mult_4_S5_2_inst3_MM23 inst3_net079 dp_cluster_0_mult_4_ab_3__2_ VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MMN87_dp_cluster_0_mult_4_S5_2_inst3_MM19 VSS dp_cluster_0_mult_4_ab_2__3_ inst3_net067 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN88_dp_cluster_0_mult_4_S5_2_inst3_MM18 VSS n30 inst3_net067 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN89_dp_cluster_0_mult_4_S5_2_inst3_MM17 VSS dp_cluster_0_mult_4_ab_3__2_ inst3_net067 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN90_dp_cluster_0_mult_4_S5_2_inst3_MM16 inst3_net067 n46 n45 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN91_dp_cluster_0_mult_4_S5_2_inst3_MM11 VSS n30 inst3_net25 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN92_dp_cluster_0_mult_4_S5_2_inst3_MM10 VSS n30 inst3_net36 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN93_dp_cluster_0_mult_4_S5_2_inst3_MM9 VSS dp_cluster_0_mult_4_ab_3__2_ inst3_net25 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN94_dp_cluster_0_mult_4_S5_2_inst3_MM8 inst3_net36 dp_cluster_0_mult_4_ab_3__2_ n46 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN95_dp_cluster_0_mult_4_S5_2_inst3_MM7 inst3_net25 dp_cluster_0_mult_4_ab_2__3_ n46 VSS nmos_lvt w=54.0n l=20n nfin=2

* FAxp33_ASAP7_6t_L dp_cluster_0_mult_4_S4_1
MMP96_dp_cluster_0_mult_4_S4_1_inst4_MM22 n47 n31 inst4_net081 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP97_dp_cluster_0_mult_4_S4_1_inst4_MM21 inst4_net081 n28 inst4_net082 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP98_dp_cluster_0_mult_4_S4_1_inst4_MM20 inst4_net082 dp_cluster_0_mult_4_ab_3__1_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP99_dp_cluster_0_mult_4_S4_1_inst4_MM15 n47 n48 inst4_net027 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP100_dp_cluster_0_mult_4_S4_1_inst4_MM14 inst4_net027 n31 VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP101_dp_cluster_0_mult_4_S4_1_inst4_MM13 inst4_net027 n28 VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP102_dp_cluster_0_mult_4_S4_1_inst4_MM12 inst4_net027 dp_cluster_0_mult_4_ab_3__1_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP103_dp_cluster_0_mult_4_S4_1_inst4_MM5 n48 dp_cluster_0_mult_4_ab_3__1_ inst4_net37 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP104_dp_cluster_0_mult_4_S4_1_inst4_MM6 inst4_net37 n28 VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP105_dp_cluster_0_mult_4_S4_1_inst4_MM2 inst4_net27 n28 VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP106_dp_cluster_0_mult_4_S4_1_inst4_MM1 n48 n31 inst4_net27 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP107_dp_cluster_0_mult_4_S4_1_inst4_MM0 inst4_net27 dp_cluster_0_mult_4_ab_3__1_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMN108_dp_cluster_0_mult_4_S4_1_inst4_MM25 n47 n31 inst4_net080 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN109_dp_cluster_0_mult_4_S4_1_inst4_MM24 inst4_net080 n28 inst4_net079 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN110_dp_cluster_0_mult_4_S4_1_inst4_MM23 inst4_net079 dp_cluster_0_mult_4_ab_3__1_ VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MMN111_dp_cluster_0_mult_4_S4_1_inst4_MM19 VSS n31 inst4_net067 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN112_dp_cluster_0_mult_4_S4_1_inst4_MM18 VSS n28 inst4_net067 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN113_dp_cluster_0_mult_4_S4_1_inst4_MM17 VSS dp_cluster_0_mult_4_ab_3__1_ inst4_net067 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN114_dp_cluster_0_mult_4_S4_1_inst4_MM16 inst4_net067 n48 n47 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN115_dp_cluster_0_mult_4_S4_1_inst4_MM11 VSS n28 inst4_net25 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN116_dp_cluster_0_mult_4_S4_1_inst4_MM10 VSS n28 inst4_net36 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN117_dp_cluster_0_mult_4_S4_1_inst4_MM9 VSS dp_cluster_0_mult_4_ab_3__1_ inst4_net25 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN118_dp_cluster_0_mult_4_S4_1_inst4_MM8 inst4_net36 dp_cluster_0_mult_4_ab_3__1_ n48 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN119_dp_cluster_0_mult_4_S4_1_inst4_MM7 inst4_net25 n31 n48 VSS nmos_lvt w=54.0n l=20n nfin=2

* FAxp33_ASAP7_6t_L dp_cluster_0_mult_4_S4_0
MMP120_dp_cluster_0_mult_4_S4_0_inst5_MM22 n49 n29 inst5_net081 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP121_dp_cluster_0_mult_4_S4_0_inst5_MM21 inst5_net081 n26 inst5_net082 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP122_dp_cluster_0_mult_4_S4_0_inst5_MM20 inst5_net082 dp_cluster_0_mult_4_ab_3__0_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP123_dp_cluster_0_mult_4_S4_0_inst5_MM15 n49 n50 inst5_net027 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP124_dp_cluster_0_mult_4_S4_0_inst5_MM14 inst5_net027 n29 VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP125_dp_cluster_0_mult_4_S4_0_inst5_MM13 inst5_net027 n26 VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP126_dp_cluster_0_mult_4_S4_0_inst5_MM12 inst5_net027 dp_cluster_0_mult_4_ab_3__0_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP127_dp_cluster_0_mult_4_S4_0_inst5_MM5 n50 dp_cluster_0_mult_4_ab_3__0_ inst5_net37 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP128_dp_cluster_0_mult_4_S4_0_inst5_MM6 inst5_net37 n26 VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP129_dp_cluster_0_mult_4_S4_0_inst5_MM2 inst5_net27 n26 VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP130_dp_cluster_0_mult_4_S4_0_inst5_MM1 n50 n29 inst5_net27 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP131_dp_cluster_0_mult_4_S4_0_inst5_MM0 inst5_net27 dp_cluster_0_mult_4_ab_3__0_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMN132_dp_cluster_0_mult_4_S4_0_inst5_MM25 n49 n29 inst5_net080 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN133_dp_cluster_0_mult_4_S4_0_inst5_MM24 inst5_net080 n26 inst5_net079 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN134_dp_cluster_0_mult_4_S4_0_inst5_MM23 inst5_net079 dp_cluster_0_mult_4_ab_3__0_ VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MMN135_dp_cluster_0_mult_4_S4_0_inst5_MM19 VSS n29 inst5_net067 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN136_dp_cluster_0_mult_4_S4_0_inst5_MM18 VSS n26 inst5_net067 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN137_dp_cluster_0_mult_4_S4_0_inst5_MM17 VSS dp_cluster_0_mult_4_ab_3__0_ inst5_net067 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN138_dp_cluster_0_mult_4_S4_0_inst5_MM16 inst5_net067 n50 n49 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN139_dp_cluster_0_mult_4_S4_0_inst5_MM11 VSS n26 inst5_net25 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN140_dp_cluster_0_mult_4_S4_0_inst5_MM10 VSS n26 inst5_net36 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN141_dp_cluster_0_mult_4_S4_0_inst5_MM9 VSS dp_cluster_0_mult_4_ab_3__0_ inst5_net25 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN142_dp_cluster_0_mult_4_S4_0_inst5_MM8 inst5_net36 dp_cluster_0_mult_4_ab_3__0_ n50 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN143_dp_cluster_0_mult_4_S4_0_inst5_MM7 inst5_net25 n29 n50 VSS nmos_lvt w=54.0n l=20n nfin=2

* AND2x2_ASAP7_6t_L U3
MMP144_U3_inst6_MM4_0 n3 inst6_net10 VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP145_U3_inst6_MM4_1 n3 inst6_net10 VDD VDD pmos_lvt w=54.00n l=20n nfin=2
MMP146_U3_inst6_MM1 inst6_net10 dp_cluster_0_mult_4_ab_0__1_ VDD VDD pmos_lvt w=27.0n l=20n nfin=1
MMP147_U3_inst6_MM0 inst6_net10 dp_cluster_0_mult_4_ab_1__0_ VDD VDD pmos_lvt w=27.0n l=20n nfin=1
MMN148_U3_inst6_MM5_0 n3 inst6_net10 VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MMN149_U3_inst6_MM5_1 n3 inst6_net10 VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MMN150_U3_inst6_MM3 inst6_net20 dp_cluster_0_mult_4_ab_1__0_ VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MMN151_U3_inst6_MM2 inst6_net10 dp_cluster_0_mult_4_ab_0__1_ inst6_net20 VSS nmos_lvt w=54.0n l=20n nfin=2

* AND2x2_ASAP7_6t_L U4
MMP152_U4_inst7_MM4_0 n4 inst7_net10 VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP153_U4_inst7_MM4_1 n4 inst7_net10 VDD VDD pmos_lvt w=54.00n l=20n nfin=2
MMP154_U4_inst7_MM1 inst7_net10 dp_cluster_0_mult_4_ab_0__2_ VDD VDD pmos_lvt w=27.0n l=20n nfin=1
MMP155_U4_inst7_MM0 inst7_net10 dp_cluster_0_mult_4_ab_1__1_ VDD VDD pmos_lvt w=27.0n l=20n nfin=1
MMN156_U4_inst7_MM5_0 n4 inst7_net10 VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MMN157_U4_inst7_MM5_1 n4 inst7_net10 VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MMN158_U4_inst7_MM3 inst7_net20 dp_cluster_0_mult_4_ab_1__1_ VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MMN159_U4_inst7_MM2 inst7_net10 dp_cluster_0_mult_4_ab_0__2_ inst7_net20 VSS nmos_lvt w=54.0n l=20n nfin=2

* XOR2xp5r_ASAP7_6t_L U5
MMP160_U5_inst8_MM4 VDD dp_cluster_0_mult_4_ab_3__3_ inst8_net019 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP161_U5_inst8_MM5 VDD n23 inst8_net019 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP162_U5_inst8_MM6 inst8_net019 inst8_net036 n5 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP163_U5_inst8_MM2 inst8_net048 n23 inst8_net036 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP164_U5_inst8_MM3 VDD dp_cluster_0_mult_4_ab_3__3_ inst8_net048 VDD pmos_lvt w=54.0n l=20n nfin=2
MMN165_U5_inst8_MM11 VSS dp_cluster_0_mult_4_ab_3__3_ inst8_net047 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN166_U5_inst8_MM10 inst8_net047 n23 n5 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN167_U5_inst8_MM9 VSS inst8_net036 n5 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN168_U5_inst8_MM0 VSS dp_cluster_0_mult_4_ab_3__3_ inst8_net036 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN169_U5_inst8_MM1 VSS n23 inst8_net036 VSS nmos_lvt w=54.0n l=20n nfin=2

* XOR2xp5r_ASAP7_6t_L U6
MMP170_U6_inst9_MM4 VDD n24 inst9_net019 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP171_U6_inst9_MM5 VDD n21 inst9_net019 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP172_U6_inst9_MM6 inst9_net019 inst9_net036 n6 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP173_U6_inst9_MM2 inst9_net048 n21 inst9_net036 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP174_U6_inst9_MM3 VDD n24 inst9_net048 VDD pmos_lvt w=54.0n l=20n nfin=2
MMN175_U6_inst9_MM11 VSS n24 inst9_net047 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN176_U6_inst9_MM10 inst9_net047 n21 n6 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN177_U6_inst9_MM9 VSS inst9_net036 n6 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN178_U6_inst9_MM0 VSS n24 inst9_net036 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN179_U6_inst9_MM1 VSS n21 inst9_net036 VSS nmos_lvt w=54.0n l=20n nfin=2

* AND2x2_ASAP7_6t_L U7
MMP180_U7_inst10_MM4_0 n7 inst10_net10 VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP181_U7_inst10_MM4_1 n7 inst10_net10 VDD VDD pmos_lvt w=54.00n l=20n nfin=2
MMP182_U7_inst10_MM1 inst10_net10 dp_cluster_0_mult_4_ab_0__3_ VDD VDD pmos_lvt w=27.0n l=20n nfin=1
MMP183_U7_inst10_MM0 inst10_net10 dp_cluster_0_mult_4_ab_1__2_ VDD VDD pmos_lvt w=27.0n l=20n nfin=1
MMN184_U7_inst10_MM5_0 n7 inst10_net10 VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MMN185_U7_inst10_MM5_1 n7 inst10_net10 VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MMN186_U7_inst10_MM3 inst10_net20 dp_cluster_0_mult_4_ab_1__2_ VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MMN187_U7_inst10_MM2 inst10_net10 dp_cluster_0_mult_4_ab_0__3_ inst10_net20 VSS nmos_lvt w=54.0n l=20n nfin=2

* XOR2xp5r_ASAP7_6t_L U8
MMP188_U8_inst11_MM4 VDD dp_cluster_0_mult_4_ab_0__2_ inst11_net019 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP189_U8_inst11_MM5 VDD dp_cluster_0_mult_4_ab_1__1_ inst11_net019 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP190_U8_inst11_MM6 inst11_net019 inst11_net036 n8 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP191_U8_inst11_MM2 inst11_net048 dp_cluster_0_mult_4_ab_1__1_ inst11_net036 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP192_U8_inst11_MM3 VDD dp_cluster_0_mult_4_ab_0__2_ inst11_net048 VDD pmos_lvt w=54.0n l=20n nfin=2
MMN193_U8_inst11_MM11 VSS dp_cluster_0_mult_4_ab_0__2_ inst11_net047 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN194_U8_inst11_MM10 inst11_net047 dp_cluster_0_mult_4_ab_1__1_ n8 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN195_U8_inst11_MM9 VSS inst11_net036 n8 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN196_U8_inst11_MM0 VSS dp_cluster_0_mult_4_ab_0__2_ inst11_net036 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN197_U8_inst11_MM1 VSS dp_cluster_0_mult_4_ab_1__1_ inst11_net036 VSS nmos_lvt w=54.0n l=20n nfin=2

* XOR2xp5r_ASAP7_6t_L U9
MMP198_U9_inst12_MM4 VDD dp_cluster_0_mult_4_ab_0__3_ inst12_net019 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP199_U9_inst12_MM5 VDD dp_cluster_0_mult_4_ab_1__2_ inst12_net019 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP200_U9_inst12_MM6 inst12_net019 inst12_net036 n9 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP201_U9_inst12_MM2 inst12_net048 dp_cluster_0_mult_4_ab_1__2_ inst12_net036 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP202_U9_inst12_MM3 VDD dp_cluster_0_mult_4_ab_0__3_ inst12_net048 VDD pmos_lvt w=54.0n l=20n nfin=2
MMN203_U9_inst12_MM11 VSS dp_cluster_0_mult_4_ab_0__3_ inst12_net047 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN204_U9_inst12_MM10 inst12_net047 dp_cluster_0_mult_4_ab_1__2_ n9 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN205_U9_inst12_MM9 VSS inst12_net036 n9 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN206_U9_inst12_MM0 VSS dp_cluster_0_mult_4_ab_0__3_ inst12_net036 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN207_U9_inst12_MM1 VSS dp_cluster_0_mult_4_ab_1__2_ inst12_net036 VSS nmos_lvt w=54.0n l=20n nfin=2

* AND2x2_ASAP7_6t_L U10
MMP208_U10_inst13_MM4_0 n10 inst13_net10 VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP209_U10_inst13_MM4_1 n10 inst13_net10 VDD VDD pmos_lvt w=54.00n l=20n nfin=2
MMP210_U10_inst13_MM1 inst13_net10 dp_cluster_0_mult_4_ab_3__3_ VDD VDD pmos_lvt w=27.0n l=20n nfin=1
MMP211_U10_inst13_MM0 inst13_net10 n23 VDD VDD pmos_lvt w=27.0n l=20n nfin=1
MMN212_U10_inst13_MM5_0 n10 inst13_net10 VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MMN213_U10_inst13_MM5_1 n10 inst13_net10 VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MMN214_U10_inst13_MM3 inst13_net20 n23 VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MMN215_U10_inst13_MM2 inst13_net10 dp_cluster_0_mult_4_ab_3__3_ inst13_net20 VSS nmos_lvt w=54.0n l=20n nfin=2

* AND2x2_ASAP7_6t_L U11
MMP216_U11_inst14_MM4_0 n11 inst14_net10 VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP217_U11_inst14_MM4_1 n11 inst14_net10 VDD VDD pmos_lvt w=54.00n l=20n nfin=2
MMP218_U11_inst14_MM1 inst14_net10 n24 VDD VDD pmos_lvt w=27.0n l=20n nfin=1
MMP219_U11_inst14_MM0 inst14_net10 n21 VDD VDD pmos_lvt w=27.0n l=20n nfin=1
MMN220_U11_inst14_MM5_0 n11 inst14_net10 VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MMN221_U11_inst14_MM5_1 n11 inst14_net10 VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MMN222_U11_inst14_MM3 inst14_net20 n21 VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MMN223_U11_inst14_MM2 inst14_net10 n24 inst14_net20 VSS nmos_lvt w=54.0n l=20n nfin=2

* AND2x2_ASAP7_6t_L U12
MMP224_U12_inst15_MM4_0 n12 inst15_net10 VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP225_U12_inst15_MM4_1 n12 inst15_net10 VDD VDD pmos_lvt w=54.00n l=20n nfin=2
MMP226_U12_inst15_MM1 inst15_net10 n22 VDD VDD pmos_lvt w=27.0n l=20n nfin=1
MMP227_U12_inst15_MM0 inst15_net10 n18 VDD VDD pmos_lvt w=27.0n l=20n nfin=1
MMN228_U12_inst15_MM5_0 n12 inst15_net10 VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MMN229_U12_inst15_MM5_1 n12 inst15_net10 VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MMN230_U12_inst15_MM3 inst15_net20 n18 VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MMN231_U12_inst15_MM2 inst15_net10 n22 inst15_net20 VSS nmos_lvt w=54.0n l=20n nfin=2

* OR2x2_ASAP7_6t_L U13
MMN232_U13_inst16_MM5_1 VSS inst16_net7 n13 VSS nmos_lvt w=54.00n l=20n nfin=2
MMN233_U13_inst16_MM5_2 VSS inst16_net7 n13 VSS nmos_lvt w=54.00n l=20n nfin=2
MMN234_U13_inst16_MM1 VSS n6 inst16_net7 VSS nmos_lvt w=27.0n l=20n nfin=1
MMN235_U13_inst16_MM2 VSS n12 inst16_net7 VSS nmos_lvt w=27.0n l=20n nfin=1
MMP236_U13_inst16_MM0_1 VDD inst16_net7 n13 VDD pmos_lvt w=54.00n l=20n nfin=2
MMP237_U13_inst16_MM0_2 VDD inst16_net7 n13 VDD pmos_lvt w=54.00n l=20n nfin=2
MMP238_U13_inst16_MM4 inst16_net15 n6 inst16_net7 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP239_U13_inst16_MM3 VDD n12 inst16_net15 VDD pmos_lvt w=54.0n l=20n nfin=2

* XOR2xp5r_ASAP7_6t_L U14
MMP240_U14_inst17_MM4 VDD dp_cluster_0_mult_4_ab_0__1_ inst17_net019 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP241_U14_inst17_MM5 VDD dp_cluster_0_mult_4_ab_1__0_ inst17_net019 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP242_U14_inst17_MM6 inst17_net019 inst17_net036 y_1_ VDD pmos_lvt w=54.0n l=20n nfin=2
MMP243_U14_inst17_MM2 inst17_net048 dp_cluster_0_mult_4_ab_1__0_ inst17_net036 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP244_U14_inst17_MM3 VDD dp_cluster_0_mult_4_ab_0__1_ inst17_net048 VDD pmos_lvt w=54.0n l=20n nfin=2
MMN245_U14_inst17_MM11 VSS dp_cluster_0_mult_4_ab_0__1_ inst17_net047 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN246_U14_inst17_MM10 inst17_net047 dp_cluster_0_mult_4_ab_1__0_ y_1_ VSS nmos_lvt w=54.0n l=20n nfin=2
MMN247_U14_inst17_MM9 VSS inst17_net036 y_1_ VSS nmos_lvt w=54.0n l=20n nfin=2
MMN248_U14_inst17_MM0 VSS dp_cluster_0_mult_4_ab_0__1_ inst17_net036 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN249_U14_inst17_MM1 VSS dp_cluster_0_mult_4_ab_1__0_ inst17_net036 VSS nmos_lvt w=54.0n l=20n nfin=2

* XOR2xp5r_ASAP7_6t_L U15
MMP250_U15_inst18_MM4 VDD n22 inst18_net019 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP251_U15_inst18_MM5 VDD n18 inst18_net019 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP252_U15_inst18_MM6 inst18_net019 inst18_net036 y_4_ VDD pmos_lvt w=54.0n l=20n nfin=2
MMP253_U15_inst18_MM2 inst18_net048 n18 inst18_net036 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP254_U15_inst18_MM3 VDD n22 inst18_net048 VDD pmos_lvt w=54.0n l=20n nfin=2
MMN255_U15_inst18_MM11 VSS n22 inst18_net047 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN256_U15_inst18_MM10 inst18_net047 n18 y_4_ VSS nmos_lvt w=54.0n l=20n nfin=2
MMN257_U15_inst18_MM9 VSS inst18_net036 y_4_ VSS nmos_lvt w=54.0n l=20n nfin=2
MMN258_U15_inst18_MM0 VSS n22 inst18_net036 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN259_U15_inst18_MM1 VSS n18 inst18_net036 VSS nmos_lvt w=54.0n l=20n nfin=2

* AND2x2_ASAP7_6t_L U16
MMP260_U16_inst19_MM4_0 y_5_ inst19_net10 VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP261_U16_inst19_MM4_1 y_5_ inst19_net10 VDD VDD pmos_lvt w=54.00n l=20n nfin=2
MMP262_U16_inst19_MM1 inst19_net10 n55 VDD VDD pmos_lvt w=27.0n l=20n nfin=1
MMP263_U16_inst19_MM0 inst19_net10 n13 VDD VDD pmos_lvt w=27.0n l=20n nfin=1
MMN264_U16_inst19_MM5_0 y_5_ inst19_net10 VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MMN265_U16_inst19_MM5_1 y_5_ inst19_net10 VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MMN266_U16_inst19_MM3 inst19_net20 n13 VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MMN267_U16_inst19_MM2 inst19_net10 n55 inst19_net20 VSS nmos_lvt w=54.0n l=20n nfin=2

* OAI21xp5b_ASAP7_6t_L U17
MMP268_U17_inst20_MM2 n51 n53 VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP269_U17_inst20_MM1 n51 n55 inst20_net27 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP270_U17_inst20_MM0 inst20_net27 n52 VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMN271_U17_inst20_MM6 inst20_net11 n53 VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MMN272_U17_inst20_MM5 n51 n55 inst20_net11 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN273_U17_inst20_MM4 n51 n52 inst20_net11 VSS nmos_lvt w=54.0n l=20n nfin=2

* INVx1_ASAP7_6t_L U18
MMN274_U18_inst21_MM0 n17 n55 VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MMP275_U18_inst21_MM1 n17 n55 VDD VDD pmos_lvt w=54.0n l=20n nfin=2

* INVx1_ASAP7_6t_L U19
MMN276_U19_inst22_MM0 n18 n50 VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MMP277_U19_inst22_MM1 n18 n50 VDD VDD pmos_lvt w=54.0n l=20n nfin=2

* INVx1_ASAP7_6t_L U20
MMN278_U20_inst23_MM0 y_3_ n49 VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MMP279_U20_inst23_MM1 y_3_ n49 VDD VDD pmos_lvt w=54.0n l=20n nfin=2

* INVx1_ASAP7_6t_L U21
MMN280_U21_inst24_MM0 n20 n53 VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MMP281_U21_inst24_MM1 n20 n53 VDD VDD pmos_lvt w=54.0n l=20n nfin=2

* INVx1_ASAP7_6t_L U22
MMN282_U22_inst25_MM0 n21 n48 VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MMP283_U22_inst25_MM1 n21 n48 VDD VDD pmos_lvt w=54.0n l=20n nfin=2

* INVx1_ASAP7_6t_L U23
MMN284_U23_inst26_MM0 n22 n47 VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MMP285_U23_inst26_MM1 n22 n47 VDD VDD pmos_lvt w=54.0n l=20n nfin=2

* INVx1_ASAP7_6t_L U24
MMN286_U24_inst27_MM0 n23 n46 VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MMP287_U24_inst27_MM1 n23 n46 VDD VDD pmos_lvt w=54.0n l=20n nfin=2

* INVx1_ASAP7_6t_L U25
MMN288_U25_inst28_MM0 n24 n45 VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MMP289_U25_inst28_MM1 n24 n45 VDD VDD pmos_lvt w=54.0n l=20n nfin=2

* INVx1_ASAP7_6t_L U26
MMN290_U26_inst29_MM0 n25 a_3_ VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MMP291_U26_inst29_MM1 n25 a_3_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2

* INVx1_ASAP7_6t_L U27
MMN292_U27_inst30_MM0 n26 n44 VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MMP293_U27_inst30_MM1 n26 n44 VDD VDD pmos_lvt w=54.0n l=20n nfin=2

* INVx1_ASAP7_6t_L U28
MMN294_U28_inst31_MM0 y_2_ n43 VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MMP295_U28_inst31_MM1 y_2_ n43 VDD VDD pmos_lvt w=54.0n l=20n nfin=2

* INVx1_ASAP7_6t_L U29
MMN296_U29_inst32_MM0 n28 n42 VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MMP297_U29_inst32_MM1 n28 n42 VDD VDD pmos_lvt w=54.0n l=20n nfin=2

* INVx1_ASAP7_6t_L U30
MMN298_U30_inst33_MM0 n29 n41 VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MMP299_U30_inst33_MM1 n29 n41 VDD VDD pmos_lvt w=54.0n l=20n nfin=2

* INVx1_ASAP7_6t_L U31
MMN300_U31_inst34_MM0 n30 n40 VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MMP301_U31_inst34_MM1 n30 n40 VDD VDD pmos_lvt w=54.0n l=20n nfin=2

* INVx1_ASAP7_6t_L U32
MMN302_U32_inst35_MM0 n31 n39 VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MMP303_U32_inst35_MM1 n31 n39 VDD VDD pmos_lvt w=54.0n l=20n nfin=2

* INVx1_ASAP7_6t_L U33
MMN304_U33_inst36_MM0 n32 a_2_ VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MMP305_U33_inst36_MM1 n32 a_2_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2

* INVx1_ASAP7_6t_L U34
MMN306_U34_inst37_MM0 n33 a_1_ VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MMP307_U34_inst37_MM1 n33 a_1_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2

* INVx1_ASAP7_6t_L U35
MMN308_U35_inst38_MM0 n34 a_0_ VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MMP309_U35_inst38_MM1 n34 a_0_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2

* INVx1_ASAP7_6t_L U36
MMN310_U36_inst39_MM0 n35 b_3_ VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MMP311_U36_inst39_MM1 n35 b_3_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2

* INVx1_ASAP7_6t_L U37
MMN312_U37_inst40_MM0 n36 b_2_ VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MMP313_U37_inst40_MM1 n36 b_2_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2

* INVx1_ASAP7_6t_L U38
MMN314_U38_inst41_MM0 n37 b_1_ VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MMP315_U38_inst41_MM1 n37 b_1_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2

* INVx1_ASAP7_6t_L U39
MMN316_U39_inst42_MM0 n38 b_0_ VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MMP317_U39_inst42_MM1 n38 b_0_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2

* NOR2xp5_ASAP7_6t_L U40
MMN318_U40_inst43_MM2 VSS n38 y_0_ VSS nmos_lvt w=27.0n l=20n nfin=1
MMN319_U40_inst43_MM1 VSS n34 y_0_ VSS nmos_lvt w=27.0n l=20n nfin=1
MMP320_U40_inst43_MM4 inst43_net16 n34 y_0_ VDD pmos_lvt w=54.0n l=20n nfin=2
MMP321_U40_inst43_MM3 VDD n38 inst43_net16 VDD pmos_lvt w=54.0n l=20n nfin=2

* NOR2xp5_ASAP7_6t_L U41
MMN322_U41_inst44_MM2 VSS n37 dp_cluster_0_mult_4_ab_0__1_ VSS nmos_lvt w=27.0n l=20n nfin=1
MMN323_U41_inst44_MM1 VSS n34 dp_cluster_0_mult_4_ab_0__1_ VSS nmos_lvt w=27.0n l=20n nfin=1
MMP324_U41_inst44_MM4 inst44_net16 n34 dp_cluster_0_mult_4_ab_0__1_ VDD pmos_lvt w=54.0n l=20n nfin=2
MMP325_U41_inst44_MM3 VDD n37 inst44_net16 VDD pmos_lvt w=54.0n l=20n nfin=2

* NOR2xp5_ASAP7_6t_L U42
MMN326_U42_inst45_MM2 VSS n36 dp_cluster_0_mult_4_ab_0__2_ VSS nmos_lvt w=27.0n l=20n nfin=1
MMN327_U42_inst45_MM1 VSS n34 dp_cluster_0_mult_4_ab_0__2_ VSS nmos_lvt w=27.0n l=20n nfin=1
MMP328_U42_inst45_MM4 inst45_net16 n34 dp_cluster_0_mult_4_ab_0__2_ VDD pmos_lvt w=54.0n l=20n nfin=2
MMP329_U42_inst45_MM3 VDD n36 inst45_net16 VDD pmos_lvt w=54.0n l=20n nfin=2

* NOR2xp5_ASAP7_6t_L U43
MMN330_U43_inst46_MM2 VSS n35 dp_cluster_0_mult_4_ab_0__3_ VSS nmos_lvt w=27.0n l=20n nfin=1
MMN331_U43_inst46_MM1 VSS n34 dp_cluster_0_mult_4_ab_0__3_ VSS nmos_lvt w=27.0n l=20n nfin=1
MMP332_U43_inst46_MM4 inst46_net16 n34 dp_cluster_0_mult_4_ab_0__3_ VDD pmos_lvt w=54.0n l=20n nfin=2
MMP333_U43_inst46_MM3 VDD n35 inst46_net16 VDD pmos_lvt w=54.0n l=20n nfin=2

* NOR2xp5_ASAP7_6t_L U44
MMN334_U44_inst47_MM2 VSS n38 dp_cluster_0_mult_4_ab_1__0_ VSS nmos_lvt w=27.0n l=20n nfin=1
MMN335_U44_inst47_MM1 VSS n33 dp_cluster_0_mult_4_ab_1__0_ VSS nmos_lvt w=27.0n l=20n nfin=1
MMP336_U44_inst47_MM4 inst47_net16 n33 dp_cluster_0_mult_4_ab_1__0_ VDD pmos_lvt w=54.0n l=20n nfin=2
MMP337_U44_inst47_MM3 VDD n38 inst47_net16 VDD pmos_lvt w=54.0n l=20n nfin=2

* NOR2xp5_ASAP7_6t_L U45
MMN338_U45_inst48_MM2 VSS n37 dp_cluster_0_mult_4_ab_1__1_ VSS nmos_lvt w=27.0n l=20n nfin=1
MMN339_U45_inst48_MM1 VSS n33 dp_cluster_0_mult_4_ab_1__1_ VSS nmos_lvt w=27.0n l=20n nfin=1
MMP340_U45_inst48_MM4 inst48_net16 n33 dp_cluster_0_mult_4_ab_1__1_ VDD pmos_lvt w=54.0n l=20n nfin=2
MMP341_U45_inst48_MM3 VDD n37 inst48_net16 VDD pmos_lvt w=54.0n l=20n nfin=2

* NOR2xp5_ASAP7_6t_L U46
MMN342_U46_inst49_MM2 VSS n36 dp_cluster_0_mult_4_ab_1__2_ VSS nmos_lvt w=27.0n l=20n nfin=1
MMN343_U46_inst49_MM1 VSS n33 dp_cluster_0_mult_4_ab_1__2_ VSS nmos_lvt w=27.0n l=20n nfin=1
MMP344_U46_inst49_MM4 inst49_net16 n33 dp_cluster_0_mult_4_ab_1__2_ VDD pmos_lvt w=54.0n l=20n nfin=2
MMP345_U46_inst49_MM3 VDD n36 inst49_net16 VDD pmos_lvt w=54.0n l=20n nfin=2

* NOR2xp5_ASAP7_6t_L U47
MMN346_U47_inst50_MM2 VSS n35 dp_cluster_0_mult_4_ab_1__3_ VSS nmos_lvt w=27.0n l=20n nfin=1
MMN347_U47_inst50_MM1 VSS n33 dp_cluster_0_mult_4_ab_1__3_ VSS nmos_lvt w=27.0n l=20n nfin=1
MMP348_U47_inst50_MM4 inst50_net16 n33 dp_cluster_0_mult_4_ab_1__3_ VDD pmos_lvt w=54.0n l=20n nfin=2
MMP349_U47_inst50_MM3 VDD n35 inst50_net16 VDD pmos_lvt w=54.0n l=20n nfin=2

* NOR2xp5_ASAP7_6t_L U48
MMN350_U48_inst51_MM2 VSS n38 dp_cluster_0_mult_4_ab_2__0_ VSS nmos_lvt w=27.0n l=20n nfin=1
MMN351_U48_inst51_MM1 VSS n32 dp_cluster_0_mult_4_ab_2__0_ VSS nmos_lvt w=27.0n l=20n nfin=1
MMP352_U48_inst51_MM4 inst51_net16 n32 dp_cluster_0_mult_4_ab_2__0_ VDD pmos_lvt w=54.0n l=20n nfin=2
MMP353_U48_inst51_MM3 VDD n38 inst51_net16 VDD pmos_lvt w=54.0n l=20n nfin=2

* NOR2xp5_ASAP7_6t_L U49
MMN354_U49_inst52_MM2 VSS n37 dp_cluster_0_mult_4_ab_2__1_ VSS nmos_lvt w=27.0n l=20n nfin=1
MMN355_U49_inst52_MM1 VSS n32 dp_cluster_0_mult_4_ab_2__1_ VSS nmos_lvt w=27.0n l=20n nfin=1
MMP356_U49_inst52_MM4 inst52_net16 n32 dp_cluster_0_mult_4_ab_2__1_ VDD pmos_lvt w=54.0n l=20n nfin=2
MMP357_U49_inst52_MM3 VDD n37 inst52_net16 VDD pmos_lvt w=54.0n l=20n nfin=2

* NOR2xp5_ASAP7_6t_L U50
MMN358_U50_inst53_MM2 VSS n36 dp_cluster_0_mult_4_ab_2__2_ VSS nmos_lvt w=27.0n l=20n nfin=1
MMN359_U50_inst53_MM1 VSS n32 dp_cluster_0_mult_4_ab_2__2_ VSS nmos_lvt w=27.0n l=20n nfin=1
MMP360_U50_inst53_MM4 inst53_net16 n32 dp_cluster_0_mult_4_ab_2__2_ VDD pmos_lvt w=54.0n l=20n nfin=2
MMP361_U50_inst53_MM3 VDD n36 inst53_net16 VDD pmos_lvt w=54.0n l=20n nfin=2

* NOR2xp5_ASAP7_6t_L U51
MMN362_U51_inst54_MM2 VSS n35 dp_cluster_0_mult_4_ab_2__3_ VSS nmos_lvt w=27.0n l=20n nfin=1
MMN363_U51_inst54_MM1 VSS n32 dp_cluster_0_mult_4_ab_2__3_ VSS nmos_lvt w=27.0n l=20n nfin=1
MMP364_U51_inst54_MM4 inst54_net16 n32 dp_cluster_0_mult_4_ab_2__3_ VDD pmos_lvt w=54.0n l=20n nfin=2
MMP365_U51_inst54_MM3 VDD n35 inst54_net16 VDD pmos_lvt w=54.0n l=20n nfin=2

* NOR2xp5_ASAP7_6t_L U52
MMN366_U52_inst55_MM2 VSS n25 dp_cluster_0_mult_4_ab_3__0_ VSS nmos_lvt w=27.0n l=20n nfin=1
MMN367_U52_inst55_MM1 VSS n38 dp_cluster_0_mult_4_ab_3__0_ VSS nmos_lvt w=27.0n l=20n nfin=1
MMP368_U52_inst55_MM4 inst55_net16 n38 dp_cluster_0_mult_4_ab_3__0_ VDD pmos_lvt w=54.0n l=20n nfin=2
MMP369_U52_inst55_MM3 VDD n25 inst55_net16 VDD pmos_lvt w=54.0n l=20n nfin=2

* NOR2xp5_ASAP7_6t_L U53
MMN370_U53_inst56_MM2 VSS n25 dp_cluster_0_mult_4_ab_3__1_ VSS nmos_lvt w=27.0n l=20n nfin=1
MMN371_U53_inst56_MM1 VSS n37 dp_cluster_0_mult_4_ab_3__1_ VSS nmos_lvt w=27.0n l=20n nfin=1
MMP372_U53_inst56_MM4 inst56_net16 n37 dp_cluster_0_mult_4_ab_3__1_ VDD pmos_lvt w=54.0n l=20n nfin=2
MMP373_U53_inst56_MM3 VDD n25 inst56_net16 VDD pmos_lvt w=54.0n l=20n nfin=2

* NOR2xp5_ASAP7_6t_L U54
MMN374_U54_inst57_MM2 VSS n25 dp_cluster_0_mult_4_ab_3__2_ VSS nmos_lvt w=27.0n l=20n nfin=1
MMN375_U54_inst57_MM1 VSS n36 dp_cluster_0_mult_4_ab_3__2_ VSS nmos_lvt w=27.0n l=20n nfin=1
MMP376_U54_inst57_MM4 inst57_net16 n36 dp_cluster_0_mult_4_ab_3__2_ VDD pmos_lvt w=54.0n l=20n nfin=2
MMP377_U54_inst57_MM3 VDD n25 inst57_net16 VDD pmos_lvt w=54.0n l=20n nfin=2

* NOR2xp5_ASAP7_6t_L U55
MMN378_U55_inst58_MM2 VSS n25 dp_cluster_0_mult_4_ab_3__3_ VSS nmos_lvt w=27.0n l=20n nfin=1
MMN379_U55_inst58_MM1 VSS n35 dp_cluster_0_mult_4_ab_3__3_ VSS nmos_lvt w=27.0n l=20n nfin=1
MMP380_U55_inst58_MM4 inst58_net16 n35 dp_cluster_0_mult_4_ab_3__3_ VDD pmos_lvt w=54.0n l=20n nfin=2
MMP381_U55_inst58_MM3 VDD n25 inst58_net16 VDD pmos_lvt w=54.0n l=20n nfin=2

* XOR2xp5r_ASAP7_6t_L U56
MMP382_U56_inst59_MM4 VDD n10 inst59_net019 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP383_U56_inst59_MM5 VDD n51 inst59_net019 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP384_U56_inst59_MM6 inst59_net019 inst59_net036 y_7_ VDD pmos_lvt w=54.0n l=20n nfin=2
MMP385_U56_inst59_MM2 inst59_net048 n51 inst59_net036 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP386_U56_inst59_MM3 VDD n10 inst59_net048 VDD pmos_lvt w=54.0n l=20n nfin=2
MMN387_U56_inst59_MM11 VSS n10 inst59_net047 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN388_U56_inst59_MM10 inst59_net047 n51 y_7_ VSS nmos_lvt w=54.0n l=20n nfin=2
MMN389_U56_inst59_MM9 VSS inst59_net036 y_7_ VSS nmos_lvt w=54.0n l=20n nfin=2
MMN390_U56_inst59_MM0 VSS n10 inst59_net036 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN391_U56_inst59_MM1 VSS n51 inst59_net036 VSS nmos_lvt w=54.0n l=20n nfin=2

* XOR2xp5r_ASAP7_6t_L U57
MMP392_U57_inst60_MM4 VDD n54 inst60_net019 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP393_U57_inst60_MM5 VDD n17 inst60_net019 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP394_U57_inst60_MM6 inst60_net019 inst60_net036 y_6_ VDD pmos_lvt w=54.0n l=20n nfin=2
MMP395_U57_inst60_MM2 inst60_net048 n17 inst60_net036 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP396_U57_inst60_MM3 VDD n54 inst60_net048 VDD pmos_lvt w=54.0n l=20n nfin=2
MMN397_U57_inst60_MM11 VSS n54 inst60_net047 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN398_U57_inst60_MM10 inst60_net047 n17 y_6_ VSS nmos_lvt w=54.0n l=20n nfin=2
MMN399_U57_inst60_MM9 VSS inst60_net036 y_6_ VSS nmos_lvt w=54.0n l=20n nfin=2
MMN400_U57_inst60_MM0 VSS n54 inst60_net036 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN401_U57_inst60_MM1 VSS n17 inst60_net036 VSS nmos_lvt w=54.0n l=20n nfin=2

* NOR2xp5_ASAP7_6t_L U58
MMN402_U58_inst61_MM2 VSS n20 n54 VSS nmos_lvt w=27.0n l=20n nfin=1
MMN403_U58_inst61_MM1 VSS n52 n54 VSS nmos_lvt w=27.0n l=20n nfin=1
MMP404_U58_inst61_MM4 inst61_net16 n52 n54 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP405_U58_inst61_MM3 VDD n20 inst61_net16 VDD pmos_lvt w=54.0n l=20n nfin=2

* NOR2xp5_ASAP7_6t_L U59
MMN406_U59_inst62_MM2 VSS n11 n52 VSS nmos_lvt w=27.0n l=20n nfin=1
MMN407_U59_inst62_MM1 VSS n5 n52 VSS nmos_lvt w=27.0n l=20n nfin=1
MMP408_U59_inst62_MM4 inst62_net16 n5 n52 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP409_U59_inst62_MM3 VDD n11 inst62_net16 VDD pmos_lvt w=54.0n l=20n nfin=2

* NAND2xp5R_ASAP7_6t_L U60
MMN410_U60_inst63_MM3 inst63_net16 n11 VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MMN411_U60_inst63_MM2 n53 n5 inst63_net16 VSS nmos_lvt w=54.0n l=20n nfin=2
MMP412_U60_inst63_MM1 n53 n5 VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP413_U60_inst63_MM0 n53 n11 VDD VDD pmos_lvt w=54.0n l=20n nfin=2

* NAND2xp5R_ASAP7_6t_L U61
MMN414_U61_inst64_MM3 inst64_net16 n12 VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MMN415_U61_inst64_MM2 n55 n6 inst64_net16 VSS nmos_lvt w=54.0n l=20n nfin=2
MMP416_U61_inst64_MM1 n55 n6 VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP417_U61_inst64_MM0 n55 n12 VDD VDD pmos_lvt w=54.0n l=20n nfin=2

.ENDS
