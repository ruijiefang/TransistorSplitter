.SUBCKT adder16 a_15_ a_14_ a_13_ a_12_ a_11_ a_10_ a_9_ a_8_ a_7_ a_6_ a_5_ a_4_ a_3_ a_2_ a_1_ a_0_ b_15_ b_14_ b_13_ b_12_ b_11_ b_10_ b_9_ b_8_ b_7_ b_6_ b_5_ b_4_ b_3_ b_2_ b_1_ b_0_ y_15_ y_14_ y_13_ y_12_ y_11_ y_10_ y_9_ y_8_ y_7_ y_6_ y_5_ y_4_ y_3_ y_2_ y_1_ y_0_


* FAxp33_ASAP7_6t_L add_4_U1_0
MMP0_add_4_U1_0_inst0_MM22 n34 add_4_CI inst0_net081 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP1_add_4_U1_0_inst0_MM21 inst0_net081 b_0_ inst0_net082 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP2_add_4_U1_0_inst0_MM20 inst0_net082 a_0_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP3_add_4_U1_0_inst0_MM15 n34 n35 inst0_net027 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP4_add_4_U1_0_inst0_MM14 inst0_net027 add_4_CI VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP5_add_4_U1_0_inst0_MM13 inst0_net027 b_0_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP6_add_4_U1_0_inst0_MM12 inst0_net027 a_0_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP7_add_4_U1_0_inst0_MM5 n35 a_0_ inst0_net37 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP8_add_4_U1_0_inst0_MM6 inst0_net37 b_0_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP9_add_4_U1_0_inst0_MM2 inst0_net27 b_0_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP10_add_4_U1_0_inst0_MM1 n35 add_4_CI inst0_net27 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP11_add_4_U1_0_inst0_MM0 inst0_net27 a_0_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMN12_add_4_U1_0_inst0_MM25 n34 add_4_CI inst0_net080 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN13_add_4_U1_0_inst0_MM24 inst0_net080 b_0_ inst0_net079 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN14_add_4_U1_0_inst0_MM23 inst0_net079 a_0_ VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MMN15_add_4_U1_0_inst0_MM19 VSS add_4_CI inst0_net067 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN16_add_4_U1_0_inst0_MM18 VSS b_0_ inst0_net067 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN17_add_4_U1_0_inst0_MM17 VSS a_0_ inst0_net067 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN18_add_4_U1_0_inst0_MM16 inst0_net067 n35 n34 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN19_add_4_U1_0_inst0_MM11 VSS b_0_ inst0_net25 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN20_add_4_U1_0_inst0_MM10 VSS b_0_ inst0_net36 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN21_add_4_U1_0_inst0_MM9 VSS a_0_ inst0_net25 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN22_add_4_U1_0_inst0_MM8 inst0_net36 a_0_ n35 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN23_add_4_U1_0_inst0_MM7 inst0_net25 add_4_CI n35 VSS nmos_lvt w=54.0n l=20n nfin=2

* FAxp33_ASAP7_6t_L add_4_U1_1
MMP24_add_4_U1_1_inst1_MM22 n36 n32 inst1_net081 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP25_add_4_U1_1_inst1_MM21 inst1_net081 b_1_ inst1_net082 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP26_add_4_U1_1_inst1_MM20 inst1_net082 a_1_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP27_add_4_U1_1_inst1_MM15 n36 n37 inst1_net027 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP28_add_4_U1_1_inst1_MM14 inst1_net027 n32 VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP29_add_4_U1_1_inst1_MM13 inst1_net027 b_1_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP30_add_4_U1_1_inst1_MM12 inst1_net027 a_1_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP31_add_4_U1_1_inst1_MM5 n37 a_1_ inst1_net37 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP32_add_4_U1_1_inst1_MM6 inst1_net37 b_1_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP33_add_4_U1_1_inst1_MM2 inst1_net27 b_1_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP34_add_4_U1_1_inst1_MM1 n37 n32 inst1_net27 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP35_add_4_U1_1_inst1_MM0 inst1_net27 a_1_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMN36_add_4_U1_1_inst1_MM25 n36 n32 inst1_net080 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN37_add_4_U1_1_inst1_MM24 inst1_net080 b_1_ inst1_net079 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN38_add_4_U1_1_inst1_MM23 inst1_net079 a_1_ VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MMN39_add_4_U1_1_inst1_MM19 VSS n32 inst1_net067 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN40_add_4_U1_1_inst1_MM18 VSS b_1_ inst1_net067 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN41_add_4_U1_1_inst1_MM17 VSS a_1_ inst1_net067 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN42_add_4_U1_1_inst1_MM16 inst1_net067 n37 n36 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN43_add_4_U1_1_inst1_MM11 VSS b_1_ inst1_net25 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN44_add_4_U1_1_inst1_MM10 VSS b_1_ inst1_net36 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN45_add_4_U1_1_inst1_MM9 VSS a_1_ inst1_net25 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN46_add_4_U1_1_inst1_MM8 inst1_net36 a_1_ n37 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN47_add_4_U1_1_inst1_MM7 inst1_net25 n32 n37 VSS nmos_lvt w=54.0n l=20n nfin=2

* FAxp33_ASAP7_6t_L add_4_U1_2
MMP48_add_4_U1_2_inst2_MM22 n38 n30 inst2_net081 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP49_add_4_U1_2_inst2_MM21 inst2_net081 b_2_ inst2_net082 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP50_add_4_U1_2_inst2_MM20 inst2_net082 a_2_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP51_add_4_U1_2_inst2_MM15 n38 n39 inst2_net027 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP52_add_4_U1_2_inst2_MM14 inst2_net027 n30 VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP53_add_4_U1_2_inst2_MM13 inst2_net027 b_2_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP54_add_4_U1_2_inst2_MM12 inst2_net027 a_2_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP55_add_4_U1_2_inst2_MM5 n39 a_2_ inst2_net37 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP56_add_4_U1_2_inst2_MM6 inst2_net37 b_2_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP57_add_4_U1_2_inst2_MM2 inst2_net27 b_2_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP58_add_4_U1_2_inst2_MM1 n39 n30 inst2_net27 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP59_add_4_U1_2_inst2_MM0 inst2_net27 a_2_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMN60_add_4_U1_2_inst2_MM25 n38 n30 inst2_net080 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN61_add_4_U1_2_inst2_MM24 inst2_net080 b_2_ inst2_net079 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN62_add_4_U1_2_inst2_MM23 inst2_net079 a_2_ VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MMN63_add_4_U1_2_inst2_MM19 VSS n30 inst2_net067 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN64_add_4_U1_2_inst2_MM18 VSS b_2_ inst2_net067 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN65_add_4_U1_2_inst2_MM17 VSS a_2_ inst2_net067 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN66_add_4_U1_2_inst2_MM16 inst2_net067 n39 n38 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN67_add_4_U1_2_inst2_MM11 VSS b_2_ inst2_net25 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN68_add_4_U1_2_inst2_MM10 VSS b_2_ inst2_net36 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN69_add_4_U1_2_inst2_MM9 VSS a_2_ inst2_net25 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN70_add_4_U1_2_inst2_MM8 inst2_net36 a_2_ n39 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN71_add_4_U1_2_inst2_MM7 inst2_net25 n30 n39 VSS nmos_lvt w=54.0n l=20n nfin=2

* FAxp33_ASAP7_6t_L add_4_U1_3
MMP72_add_4_U1_3_inst3_MM22 n40 n28 inst3_net081 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP73_add_4_U1_3_inst3_MM21 inst3_net081 b_3_ inst3_net082 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP74_add_4_U1_3_inst3_MM20 inst3_net082 a_3_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP75_add_4_U1_3_inst3_MM15 n40 n41 inst3_net027 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP76_add_4_U1_3_inst3_MM14 inst3_net027 n28 VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP77_add_4_U1_3_inst3_MM13 inst3_net027 b_3_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP78_add_4_U1_3_inst3_MM12 inst3_net027 a_3_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP79_add_4_U1_3_inst3_MM5 n41 a_3_ inst3_net37 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP80_add_4_U1_3_inst3_MM6 inst3_net37 b_3_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP81_add_4_U1_3_inst3_MM2 inst3_net27 b_3_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP82_add_4_U1_3_inst3_MM1 n41 n28 inst3_net27 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP83_add_4_U1_3_inst3_MM0 inst3_net27 a_3_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMN84_add_4_U1_3_inst3_MM25 n40 n28 inst3_net080 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN85_add_4_U1_3_inst3_MM24 inst3_net080 b_3_ inst3_net079 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN86_add_4_U1_3_inst3_MM23 inst3_net079 a_3_ VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MMN87_add_4_U1_3_inst3_MM19 VSS n28 inst3_net067 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN88_add_4_U1_3_inst3_MM18 VSS b_3_ inst3_net067 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN89_add_4_U1_3_inst3_MM17 VSS a_3_ inst3_net067 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN90_add_4_U1_3_inst3_MM16 inst3_net067 n41 n40 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN91_add_4_U1_3_inst3_MM11 VSS b_3_ inst3_net25 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN92_add_4_U1_3_inst3_MM10 VSS b_3_ inst3_net36 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN93_add_4_U1_3_inst3_MM9 VSS a_3_ inst3_net25 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN94_add_4_U1_3_inst3_MM8 inst3_net36 a_3_ n41 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN95_add_4_U1_3_inst3_MM7 inst3_net25 n28 n41 VSS nmos_lvt w=54.0n l=20n nfin=2

* FAxp33_ASAP7_6t_L add_4_U1_4
MMP96_add_4_U1_4_inst4_MM22 n42 n26 inst4_net081 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP97_add_4_U1_4_inst4_MM21 inst4_net081 b_4_ inst4_net082 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP98_add_4_U1_4_inst4_MM20 inst4_net082 a_4_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP99_add_4_U1_4_inst4_MM15 n42 n43 inst4_net027 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP100_add_4_U1_4_inst4_MM14 inst4_net027 n26 VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP101_add_4_U1_4_inst4_MM13 inst4_net027 b_4_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP102_add_4_U1_4_inst4_MM12 inst4_net027 a_4_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP103_add_4_U1_4_inst4_MM5 n43 a_4_ inst4_net37 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP104_add_4_U1_4_inst4_MM6 inst4_net37 b_4_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP105_add_4_U1_4_inst4_MM2 inst4_net27 b_4_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP106_add_4_U1_4_inst4_MM1 n43 n26 inst4_net27 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP107_add_4_U1_4_inst4_MM0 inst4_net27 a_4_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMN108_add_4_U1_4_inst4_MM25 n42 n26 inst4_net080 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN109_add_4_U1_4_inst4_MM24 inst4_net080 b_4_ inst4_net079 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN110_add_4_U1_4_inst4_MM23 inst4_net079 a_4_ VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MMN111_add_4_U1_4_inst4_MM19 VSS n26 inst4_net067 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN112_add_4_U1_4_inst4_MM18 VSS b_4_ inst4_net067 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN113_add_4_U1_4_inst4_MM17 VSS a_4_ inst4_net067 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN114_add_4_U1_4_inst4_MM16 inst4_net067 n43 n42 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN115_add_4_U1_4_inst4_MM11 VSS b_4_ inst4_net25 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN116_add_4_U1_4_inst4_MM10 VSS b_4_ inst4_net36 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN117_add_4_U1_4_inst4_MM9 VSS a_4_ inst4_net25 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN118_add_4_U1_4_inst4_MM8 inst4_net36 a_4_ n43 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN119_add_4_U1_4_inst4_MM7 inst4_net25 n26 n43 VSS nmos_lvt w=54.0n l=20n nfin=2

* FAxp33_ASAP7_6t_L add_4_U1_5
MMP120_add_4_U1_5_inst5_MM22 n44 n24 inst5_net081 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP121_add_4_U1_5_inst5_MM21 inst5_net081 b_5_ inst5_net082 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP122_add_4_U1_5_inst5_MM20 inst5_net082 a_5_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP123_add_4_U1_5_inst5_MM15 n44 n45 inst5_net027 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP124_add_4_U1_5_inst5_MM14 inst5_net027 n24 VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP125_add_4_U1_5_inst5_MM13 inst5_net027 b_5_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP126_add_4_U1_5_inst5_MM12 inst5_net027 a_5_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP127_add_4_U1_5_inst5_MM5 n45 a_5_ inst5_net37 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP128_add_4_U1_5_inst5_MM6 inst5_net37 b_5_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP129_add_4_U1_5_inst5_MM2 inst5_net27 b_5_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP130_add_4_U1_5_inst5_MM1 n45 n24 inst5_net27 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP131_add_4_U1_5_inst5_MM0 inst5_net27 a_5_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMN132_add_4_U1_5_inst5_MM25 n44 n24 inst5_net080 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN133_add_4_U1_5_inst5_MM24 inst5_net080 b_5_ inst5_net079 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN134_add_4_U1_5_inst5_MM23 inst5_net079 a_5_ VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MMN135_add_4_U1_5_inst5_MM19 VSS n24 inst5_net067 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN136_add_4_U1_5_inst5_MM18 VSS b_5_ inst5_net067 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN137_add_4_U1_5_inst5_MM17 VSS a_5_ inst5_net067 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN138_add_4_U1_5_inst5_MM16 inst5_net067 n45 n44 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN139_add_4_U1_5_inst5_MM11 VSS b_5_ inst5_net25 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN140_add_4_U1_5_inst5_MM10 VSS b_5_ inst5_net36 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN141_add_4_U1_5_inst5_MM9 VSS a_5_ inst5_net25 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN142_add_4_U1_5_inst5_MM8 inst5_net36 a_5_ n45 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN143_add_4_U1_5_inst5_MM7 inst5_net25 n24 n45 VSS nmos_lvt w=54.0n l=20n nfin=2

* FAxp33_ASAP7_6t_L add_4_U1_6
MMP144_add_4_U1_6_inst6_MM22 n46 n22 inst6_net081 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP145_add_4_U1_6_inst6_MM21 inst6_net081 b_6_ inst6_net082 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP146_add_4_U1_6_inst6_MM20 inst6_net082 a_6_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP147_add_4_U1_6_inst6_MM15 n46 n47 inst6_net027 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP148_add_4_U1_6_inst6_MM14 inst6_net027 n22 VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP149_add_4_U1_6_inst6_MM13 inst6_net027 b_6_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP150_add_4_U1_6_inst6_MM12 inst6_net027 a_6_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP151_add_4_U1_6_inst6_MM5 n47 a_6_ inst6_net37 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP152_add_4_U1_6_inst6_MM6 inst6_net37 b_6_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP153_add_4_U1_6_inst6_MM2 inst6_net27 b_6_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP154_add_4_U1_6_inst6_MM1 n47 n22 inst6_net27 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP155_add_4_U1_6_inst6_MM0 inst6_net27 a_6_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMN156_add_4_U1_6_inst6_MM25 n46 n22 inst6_net080 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN157_add_4_U1_6_inst6_MM24 inst6_net080 b_6_ inst6_net079 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN158_add_4_U1_6_inst6_MM23 inst6_net079 a_6_ VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MMN159_add_4_U1_6_inst6_MM19 VSS n22 inst6_net067 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN160_add_4_U1_6_inst6_MM18 VSS b_6_ inst6_net067 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN161_add_4_U1_6_inst6_MM17 VSS a_6_ inst6_net067 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN162_add_4_U1_6_inst6_MM16 inst6_net067 n47 n46 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN163_add_4_U1_6_inst6_MM11 VSS b_6_ inst6_net25 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN164_add_4_U1_6_inst6_MM10 VSS b_6_ inst6_net36 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN165_add_4_U1_6_inst6_MM9 VSS a_6_ inst6_net25 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN166_add_4_U1_6_inst6_MM8 inst6_net36 a_6_ n47 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN167_add_4_U1_6_inst6_MM7 inst6_net25 n22 n47 VSS nmos_lvt w=54.0n l=20n nfin=2

* FAxp33_ASAP7_6t_L add_4_U1_7
MMP168_add_4_U1_7_inst7_MM22 n48 n20 inst7_net081 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP169_add_4_U1_7_inst7_MM21 inst7_net081 b_7_ inst7_net082 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP170_add_4_U1_7_inst7_MM20 inst7_net082 a_7_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP171_add_4_U1_7_inst7_MM15 n48 n49 inst7_net027 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP172_add_4_U1_7_inst7_MM14 inst7_net027 n20 VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP173_add_4_U1_7_inst7_MM13 inst7_net027 b_7_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP174_add_4_U1_7_inst7_MM12 inst7_net027 a_7_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP175_add_4_U1_7_inst7_MM5 n49 a_7_ inst7_net37 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP176_add_4_U1_7_inst7_MM6 inst7_net37 b_7_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP177_add_4_U1_7_inst7_MM2 inst7_net27 b_7_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP178_add_4_U1_7_inst7_MM1 n49 n20 inst7_net27 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP179_add_4_U1_7_inst7_MM0 inst7_net27 a_7_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMN180_add_4_U1_7_inst7_MM25 n48 n20 inst7_net080 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN181_add_4_U1_7_inst7_MM24 inst7_net080 b_7_ inst7_net079 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN182_add_4_U1_7_inst7_MM23 inst7_net079 a_7_ VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MMN183_add_4_U1_7_inst7_MM19 VSS n20 inst7_net067 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN184_add_4_U1_7_inst7_MM18 VSS b_7_ inst7_net067 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN185_add_4_U1_7_inst7_MM17 VSS a_7_ inst7_net067 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN186_add_4_U1_7_inst7_MM16 inst7_net067 n49 n48 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN187_add_4_U1_7_inst7_MM11 VSS b_7_ inst7_net25 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN188_add_4_U1_7_inst7_MM10 VSS b_7_ inst7_net36 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN189_add_4_U1_7_inst7_MM9 VSS a_7_ inst7_net25 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN190_add_4_U1_7_inst7_MM8 inst7_net36 a_7_ n49 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN191_add_4_U1_7_inst7_MM7 inst7_net25 n20 n49 VSS nmos_lvt w=54.0n l=20n nfin=2

* FAxp33_ASAP7_6t_L add_4_U1_8
MMP192_add_4_U1_8_inst8_MM22 n50 n18 inst8_net081 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP193_add_4_U1_8_inst8_MM21 inst8_net081 b_8_ inst8_net082 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP194_add_4_U1_8_inst8_MM20 inst8_net082 a_8_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP195_add_4_U1_8_inst8_MM15 n50 n51 inst8_net027 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP196_add_4_U1_8_inst8_MM14 inst8_net027 n18 VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP197_add_4_U1_8_inst8_MM13 inst8_net027 b_8_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP198_add_4_U1_8_inst8_MM12 inst8_net027 a_8_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP199_add_4_U1_8_inst8_MM5 n51 a_8_ inst8_net37 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP200_add_4_U1_8_inst8_MM6 inst8_net37 b_8_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP201_add_4_U1_8_inst8_MM2 inst8_net27 b_8_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP202_add_4_U1_8_inst8_MM1 n51 n18 inst8_net27 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP203_add_4_U1_8_inst8_MM0 inst8_net27 a_8_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMN204_add_4_U1_8_inst8_MM25 n50 n18 inst8_net080 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN205_add_4_U1_8_inst8_MM24 inst8_net080 b_8_ inst8_net079 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN206_add_4_U1_8_inst8_MM23 inst8_net079 a_8_ VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MMN207_add_4_U1_8_inst8_MM19 VSS n18 inst8_net067 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN208_add_4_U1_8_inst8_MM18 VSS b_8_ inst8_net067 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN209_add_4_U1_8_inst8_MM17 VSS a_8_ inst8_net067 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN210_add_4_U1_8_inst8_MM16 inst8_net067 n51 n50 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN211_add_4_U1_8_inst8_MM11 VSS b_8_ inst8_net25 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN212_add_4_U1_8_inst8_MM10 VSS b_8_ inst8_net36 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN213_add_4_U1_8_inst8_MM9 VSS a_8_ inst8_net25 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN214_add_4_U1_8_inst8_MM8 inst8_net36 a_8_ n51 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN215_add_4_U1_8_inst8_MM7 inst8_net25 n18 n51 VSS nmos_lvt w=54.0n l=20n nfin=2

* FAxp33_ASAP7_6t_L add_4_U1_9
MMP216_add_4_U1_9_inst9_MM22 n52 n16 inst9_net081 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP217_add_4_U1_9_inst9_MM21 inst9_net081 b_9_ inst9_net082 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP218_add_4_U1_9_inst9_MM20 inst9_net082 a_9_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP219_add_4_U1_9_inst9_MM15 n52 n53 inst9_net027 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP220_add_4_U1_9_inst9_MM14 inst9_net027 n16 VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP221_add_4_U1_9_inst9_MM13 inst9_net027 b_9_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP222_add_4_U1_9_inst9_MM12 inst9_net027 a_9_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP223_add_4_U1_9_inst9_MM5 n53 a_9_ inst9_net37 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP224_add_4_U1_9_inst9_MM6 inst9_net37 b_9_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP225_add_4_U1_9_inst9_MM2 inst9_net27 b_9_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP226_add_4_U1_9_inst9_MM1 n53 n16 inst9_net27 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP227_add_4_U1_9_inst9_MM0 inst9_net27 a_9_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMN228_add_4_U1_9_inst9_MM25 n52 n16 inst9_net080 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN229_add_4_U1_9_inst9_MM24 inst9_net080 b_9_ inst9_net079 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN230_add_4_U1_9_inst9_MM23 inst9_net079 a_9_ VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MMN231_add_4_U1_9_inst9_MM19 VSS n16 inst9_net067 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN232_add_4_U1_9_inst9_MM18 VSS b_9_ inst9_net067 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN233_add_4_U1_9_inst9_MM17 VSS a_9_ inst9_net067 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN234_add_4_U1_9_inst9_MM16 inst9_net067 n53 n52 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN235_add_4_U1_9_inst9_MM11 VSS b_9_ inst9_net25 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN236_add_4_U1_9_inst9_MM10 VSS b_9_ inst9_net36 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN237_add_4_U1_9_inst9_MM9 VSS a_9_ inst9_net25 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN238_add_4_U1_9_inst9_MM8 inst9_net36 a_9_ n53 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN239_add_4_U1_9_inst9_MM7 inst9_net25 n16 n53 VSS nmos_lvt w=54.0n l=20n nfin=2

* FAxp33_ASAP7_6t_L add_4_U1_10
MMP240_add_4_U1_10_inst10_MM22 n54 n14 inst10_net081 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP241_add_4_U1_10_inst10_MM21 inst10_net081 b_10_ inst10_net082 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP242_add_4_U1_10_inst10_MM20 inst10_net082 a_10_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP243_add_4_U1_10_inst10_MM15 n54 n55 inst10_net027 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP244_add_4_U1_10_inst10_MM14 inst10_net027 n14 VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP245_add_4_U1_10_inst10_MM13 inst10_net027 b_10_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP246_add_4_U1_10_inst10_MM12 inst10_net027 a_10_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP247_add_4_U1_10_inst10_MM5 n55 a_10_ inst10_net37 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP248_add_4_U1_10_inst10_MM6 inst10_net37 b_10_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP249_add_4_U1_10_inst10_MM2 inst10_net27 b_10_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP250_add_4_U1_10_inst10_MM1 n55 n14 inst10_net27 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP251_add_4_U1_10_inst10_MM0 inst10_net27 a_10_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMN252_add_4_U1_10_inst10_MM25 n54 n14 inst10_net080 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN253_add_4_U1_10_inst10_MM24 inst10_net080 b_10_ inst10_net079 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN254_add_4_U1_10_inst10_MM23 inst10_net079 a_10_ VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MMN255_add_4_U1_10_inst10_MM19 VSS n14 inst10_net067 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN256_add_4_U1_10_inst10_MM18 VSS b_10_ inst10_net067 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN257_add_4_U1_10_inst10_MM17 VSS a_10_ inst10_net067 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN258_add_4_U1_10_inst10_MM16 inst10_net067 n55 n54 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN259_add_4_U1_10_inst10_MM11 VSS b_10_ inst10_net25 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN260_add_4_U1_10_inst10_MM10 VSS b_10_ inst10_net36 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN261_add_4_U1_10_inst10_MM9 VSS a_10_ inst10_net25 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN262_add_4_U1_10_inst10_MM8 inst10_net36 a_10_ n55 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN263_add_4_U1_10_inst10_MM7 inst10_net25 n14 n55 VSS nmos_lvt w=54.0n l=20n nfin=2

* FAxp33_ASAP7_6t_L add_4_U1_11
MMP264_add_4_U1_11_inst11_MM22 n56 n12 inst11_net081 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP265_add_4_U1_11_inst11_MM21 inst11_net081 b_11_ inst11_net082 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP266_add_4_U1_11_inst11_MM20 inst11_net082 a_11_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP267_add_4_U1_11_inst11_MM15 n56 n57 inst11_net027 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP268_add_4_U1_11_inst11_MM14 inst11_net027 n12 VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP269_add_4_U1_11_inst11_MM13 inst11_net027 b_11_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP270_add_4_U1_11_inst11_MM12 inst11_net027 a_11_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP271_add_4_U1_11_inst11_MM5 n57 a_11_ inst11_net37 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP272_add_4_U1_11_inst11_MM6 inst11_net37 b_11_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP273_add_4_U1_11_inst11_MM2 inst11_net27 b_11_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP274_add_4_U1_11_inst11_MM1 n57 n12 inst11_net27 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP275_add_4_U1_11_inst11_MM0 inst11_net27 a_11_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMN276_add_4_U1_11_inst11_MM25 n56 n12 inst11_net080 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN277_add_4_U1_11_inst11_MM24 inst11_net080 b_11_ inst11_net079 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN278_add_4_U1_11_inst11_MM23 inst11_net079 a_11_ VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MMN279_add_4_U1_11_inst11_MM19 VSS n12 inst11_net067 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN280_add_4_U1_11_inst11_MM18 VSS b_11_ inst11_net067 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN281_add_4_U1_11_inst11_MM17 VSS a_11_ inst11_net067 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN282_add_4_U1_11_inst11_MM16 inst11_net067 n57 n56 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN283_add_4_U1_11_inst11_MM11 VSS b_11_ inst11_net25 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN284_add_4_U1_11_inst11_MM10 VSS b_11_ inst11_net36 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN285_add_4_U1_11_inst11_MM9 VSS a_11_ inst11_net25 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN286_add_4_U1_11_inst11_MM8 inst11_net36 a_11_ n57 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN287_add_4_U1_11_inst11_MM7 inst11_net25 n12 n57 VSS nmos_lvt w=54.0n l=20n nfin=2

* FAxp33_ASAP7_6t_L add_4_U1_12
MMP288_add_4_U1_12_inst12_MM22 n58 n10 inst12_net081 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP289_add_4_U1_12_inst12_MM21 inst12_net081 b_12_ inst12_net082 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP290_add_4_U1_12_inst12_MM20 inst12_net082 a_12_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP291_add_4_U1_12_inst12_MM15 n58 n59 inst12_net027 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP292_add_4_U1_12_inst12_MM14 inst12_net027 n10 VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP293_add_4_U1_12_inst12_MM13 inst12_net027 b_12_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP294_add_4_U1_12_inst12_MM12 inst12_net027 a_12_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP295_add_4_U1_12_inst12_MM5 n59 a_12_ inst12_net37 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP296_add_4_U1_12_inst12_MM6 inst12_net37 b_12_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP297_add_4_U1_12_inst12_MM2 inst12_net27 b_12_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP298_add_4_U1_12_inst12_MM1 n59 n10 inst12_net27 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP299_add_4_U1_12_inst12_MM0 inst12_net27 a_12_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMN300_add_4_U1_12_inst12_MM25 n58 n10 inst12_net080 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN301_add_4_U1_12_inst12_MM24 inst12_net080 b_12_ inst12_net079 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN302_add_4_U1_12_inst12_MM23 inst12_net079 a_12_ VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MMN303_add_4_U1_12_inst12_MM19 VSS n10 inst12_net067 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN304_add_4_U1_12_inst12_MM18 VSS b_12_ inst12_net067 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN305_add_4_U1_12_inst12_MM17 VSS a_12_ inst12_net067 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN306_add_4_U1_12_inst12_MM16 inst12_net067 n59 n58 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN307_add_4_U1_12_inst12_MM11 VSS b_12_ inst12_net25 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN308_add_4_U1_12_inst12_MM10 VSS b_12_ inst12_net36 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN309_add_4_U1_12_inst12_MM9 VSS a_12_ inst12_net25 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN310_add_4_U1_12_inst12_MM8 inst12_net36 a_12_ n59 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN311_add_4_U1_12_inst12_MM7 inst12_net25 n10 n59 VSS nmos_lvt w=54.0n l=20n nfin=2

* FAxp33_ASAP7_6t_L add_4_U1_13
MMP312_add_4_U1_13_inst13_MM22 n60 n8 inst13_net081 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP313_add_4_U1_13_inst13_MM21 inst13_net081 b_13_ inst13_net082 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP314_add_4_U1_13_inst13_MM20 inst13_net082 a_13_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP315_add_4_U1_13_inst13_MM15 n60 n61 inst13_net027 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP316_add_4_U1_13_inst13_MM14 inst13_net027 n8 VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP317_add_4_U1_13_inst13_MM13 inst13_net027 b_13_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP318_add_4_U1_13_inst13_MM12 inst13_net027 a_13_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP319_add_4_U1_13_inst13_MM5 n61 a_13_ inst13_net37 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP320_add_4_U1_13_inst13_MM6 inst13_net37 b_13_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP321_add_4_U1_13_inst13_MM2 inst13_net27 b_13_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP322_add_4_U1_13_inst13_MM1 n61 n8 inst13_net27 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP323_add_4_U1_13_inst13_MM0 inst13_net27 a_13_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMN324_add_4_U1_13_inst13_MM25 n60 n8 inst13_net080 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN325_add_4_U1_13_inst13_MM24 inst13_net080 b_13_ inst13_net079 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN326_add_4_U1_13_inst13_MM23 inst13_net079 a_13_ VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MMN327_add_4_U1_13_inst13_MM19 VSS n8 inst13_net067 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN328_add_4_U1_13_inst13_MM18 VSS b_13_ inst13_net067 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN329_add_4_U1_13_inst13_MM17 VSS a_13_ inst13_net067 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN330_add_4_U1_13_inst13_MM16 inst13_net067 n61 n60 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN331_add_4_U1_13_inst13_MM11 VSS b_13_ inst13_net25 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN332_add_4_U1_13_inst13_MM10 VSS b_13_ inst13_net36 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN333_add_4_U1_13_inst13_MM9 VSS a_13_ inst13_net25 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN334_add_4_U1_13_inst13_MM8 inst13_net36 a_13_ n61 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN335_add_4_U1_13_inst13_MM7 inst13_net25 n8 n61 VSS nmos_lvt w=54.0n l=20n nfin=2

* FAxp33_ASAP7_6t_L add_4_U1_14
MMP336_add_4_U1_14_inst14_MM22 n62 n6 inst14_net081 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP337_add_4_U1_14_inst14_MM21 inst14_net081 b_14_ inst14_net082 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP338_add_4_U1_14_inst14_MM20 inst14_net082 a_14_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP339_add_4_U1_14_inst14_MM15 n62 n63 inst14_net027 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP340_add_4_U1_14_inst14_MM14 inst14_net027 n6 VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP341_add_4_U1_14_inst14_MM13 inst14_net027 b_14_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP342_add_4_U1_14_inst14_MM12 inst14_net027 a_14_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP343_add_4_U1_14_inst14_MM5 n63 a_14_ inst14_net37 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP344_add_4_U1_14_inst14_MM6 inst14_net37 b_14_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP345_add_4_U1_14_inst14_MM2 inst14_net27 b_14_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP346_add_4_U1_14_inst14_MM1 n63 n6 inst14_net27 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP347_add_4_U1_14_inst14_MM0 inst14_net27 a_14_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMN348_add_4_U1_14_inst14_MM25 n62 n6 inst14_net080 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN349_add_4_U1_14_inst14_MM24 inst14_net080 b_14_ inst14_net079 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN350_add_4_U1_14_inst14_MM23 inst14_net079 a_14_ VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MMN351_add_4_U1_14_inst14_MM19 VSS n6 inst14_net067 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN352_add_4_U1_14_inst14_MM18 VSS b_14_ inst14_net067 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN353_add_4_U1_14_inst14_MM17 VSS a_14_ inst14_net067 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN354_add_4_U1_14_inst14_MM16 inst14_net067 n63 n62 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN355_add_4_U1_14_inst14_MM11 VSS b_14_ inst14_net25 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN356_add_4_U1_14_inst14_MM10 VSS b_14_ inst14_net36 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN357_add_4_U1_14_inst14_MM9 VSS a_14_ inst14_net25 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN358_add_4_U1_14_inst14_MM8 inst14_net36 a_14_ n63 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN359_add_4_U1_14_inst14_MM7 inst14_net25 n6 n63 VSS nmos_lvt w=54.0n l=20n nfin=2

* FAxp33_ASAP7_6t_L add_4_U1_15
MMP360_add_4_U1_15_inst15_MM22 n64 n4 inst15_net081 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP361_add_4_U1_15_inst15_MM21 inst15_net081 b_15_ inst15_net082 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP362_add_4_U1_15_inst15_MM20 inst15_net082 a_15_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP363_add_4_U1_15_inst15_MM15 n64 inst15_CON inst15_net027 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP364_add_4_U1_15_inst15_MM14 inst15_net027 n4 VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP365_add_4_U1_15_inst15_MM13 inst15_net027 b_15_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP366_add_4_U1_15_inst15_MM12 inst15_net027 a_15_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP367_add_4_U1_15_inst15_MM5 inst15_CON a_15_ inst15_net37 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP368_add_4_U1_15_inst15_MM6 inst15_net37 b_15_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP369_add_4_U1_15_inst15_MM2 inst15_net27 b_15_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMP370_add_4_U1_15_inst15_MM1 inst15_CON n4 inst15_net27 VDD pmos_lvt w=54.0n l=20n nfin=2
MMP371_add_4_U1_15_inst15_MM0 inst15_net27 a_15_ VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MMN372_add_4_U1_15_inst15_MM25 n64 n4 inst15_net080 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN373_add_4_U1_15_inst15_MM24 inst15_net080 b_15_ inst15_net079 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN374_add_4_U1_15_inst15_MM23 inst15_net079 a_15_ VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MMN375_add_4_U1_15_inst15_MM19 VSS n4 inst15_net067 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN376_add_4_U1_15_inst15_MM18 VSS b_15_ inst15_net067 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN377_add_4_U1_15_inst15_MM17 VSS a_15_ inst15_net067 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN378_add_4_U1_15_inst15_MM16 inst15_net067 inst15_CON n64 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN379_add_4_U1_15_inst15_MM11 VSS b_15_ inst15_net25 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN380_add_4_U1_15_inst15_MM10 VSS b_15_ inst15_net36 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN381_add_4_U1_15_inst15_MM9 VSS a_15_ inst15_net25 VSS nmos_lvt w=54.0n l=20n nfin=2
MMN382_add_4_U1_15_inst15_MM8 inst15_net36 a_15_ inst15_CON VSS nmos_lvt w=54.0n l=20n nfin=2
MMN383_add_4_U1_15_inst15_MM7 inst15_net25 n4 inst15_CON VSS nmos_lvt w=54.0n l=20n nfin=2

* TIELOxp5_ASAP7_6t_L U3
MMP384_U3_inst16_MM1 inst16_net9 add_4_CI VDD VDD pmos_lvt w=27.0n l=20n nfin=1
MMN385_U3_inst16_MM2 add_4_CI inst16_net9 VSS VSS nmos_lvt w=27.0n l=20n nfin=1

* INVx1_ASAP7_6t_L U4
MMN386_U4_inst17_MM0 y_15_ n64 VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MMP387_U4_inst17_MM1 y_15_ n64 VDD VDD pmos_lvt w=54.0n l=20n nfin=2

* INVx1_ASAP7_6t_L U5
MMN388_U5_inst18_MM0 n4 n63 VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MMP389_U5_inst18_MM1 n4 n63 VDD VDD pmos_lvt w=54.0n l=20n nfin=2

* INVx1_ASAP7_6t_L U6
MMN390_U6_inst19_MM0 y_14_ n62 VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MMP391_U6_inst19_MM1 y_14_ n62 VDD VDD pmos_lvt w=54.0n l=20n nfin=2

* INVx1_ASAP7_6t_L U7
MMN392_U7_inst20_MM0 n6 n61 VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MMP393_U7_inst20_MM1 n6 n61 VDD VDD pmos_lvt w=54.0n l=20n nfin=2

* INVx1_ASAP7_6t_L U8
MMN394_U8_inst21_MM0 y_13_ n60 VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MMP395_U8_inst21_MM1 y_13_ n60 VDD VDD pmos_lvt w=54.0n l=20n nfin=2

* INVx1_ASAP7_6t_L U9
MMN396_U9_inst22_MM0 n8 n59 VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MMP397_U9_inst22_MM1 n8 n59 VDD VDD pmos_lvt w=54.0n l=20n nfin=2

* INVx1_ASAP7_6t_L U10
MMN398_U10_inst23_MM0 y_12_ n58 VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MMP399_U10_inst23_MM1 y_12_ n58 VDD VDD pmos_lvt w=54.0n l=20n nfin=2

* INVx1_ASAP7_6t_L U11
MMN400_U11_inst24_MM0 n10 n57 VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MMP401_U11_inst24_MM1 n10 n57 VDD VDD pmos_lvt w=54.0n l=20n nfin=2

* INVx1_ASAP7_6t_L U12
MMN402_U12_inst25_MM0 y_11_ n56 VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MMP403_U12_inst25_MM1 y_11_ n56 VDD VDD pmos_lvt w=54.0n l=20n nfin=2

* INVx1_ASAP7_6t_L U13
MMN404_U13_inst26_MM0 n12 n55 VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MMP405_U13_inst26_MM1 n12 n55 VDD VDD pmos_lvt w=54.0n l=20n nfin=2

* INVx1_ASAP7_6t_L U14
MMN406_U14_inst27_MM0 y_10_ n54 VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MMP407_U14_inst27_MM1 y_10_ n54 VDD VDD pmos_lvt w=54.0n l=20n nfin=2

* INVx1_ASAP7_6t_L U15
MMN408_U15_inst28_MM0 n14 n53 VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MMP409_U15_inst28_MM1 n14 n53 VDD VDD pmos_lvt w=54.0n l=20n nfin=2

* INVx1_ASAP7_6t_L U16
MMN410_U16_inst29_MM0 y_9_ n52 VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MMP411_U16_inst29_MM1 y_9_ n52 VDD VDD pmos_lvt w=54.0n l=20n nfin=2

* INVx1_ASAP7_6t_L U17
MMN412_U17_inst30_MM0 n16 n51 VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MMP413_U17_inst30_MM1 n16 n51 VDD VDD pmos_lvt w=54.0n l=20n nfin=2

* INVx1_ASAP7_6t_L U18
MMN414_U18_inst31_MM0 y_8_ n50 VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MMP415_U18_inst31_MM1 y_8_ n50 VDD VDD pmos_lvt w=54.0n l=20n nfin=2

* INVx1_ASAP7_6t_L U19
MMN416_U19_inst32_MM0 n18 n49 VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MMP417_U19_inst32_MM1 n18 n49 VDD VDD pmos_lvt w=54.0n l=20n nfin=2

* INVx1_ASAP7_6t_L U20
MMN418_U20_inst33_MM0 y_7_ n48 VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MMP419_U20_inst33_MM1 y_7_ n48 VDD VDD pmos_lvt w=54.0n l=20n nfin=2

* INVx1_ASAP7_6t_L U21
MMN420_U21_inst34_MM0 n20 n47 VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MMP421_U21_inst34_MM1 n20 n47 VDD VDD pmos_lvt w=54.0n l=20n nfin=2

* INVx1_ASAP7_6t_L U22
MMN422_U22_inst35_MM0 y_6_ n46 VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MMP423_U22_inst35_MM1 y_6_ n46 VDD VDD pmos_lvt w=54.0n l=20n nfin=2

* INVx1_ASAP7_6t_L U23
MMN424_U23_inst36_MM0 n22 n45 VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MMP425_U23_inst36_MM1 n22 n45 VDD VDD pmos_lvt w=54.0n l=20n nfin=2

* INVx1_ASAP7_6t_L U24
MMN426_U24_inst37_MM0 y_5_ n44 VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MMP427_U24_inst37_MM1 y_5_ n44 VDD VDD pmos_lvt w=54.0n l=20n nfin=2

* INVx1_ASAP7_6t_L U25
MMN428_U25_inst38_MM0 n24 n43 VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MMP429_U25_inst38_MM1 n24 n43 VDD VDD pmos_lvt w=54.0n l=20n nfin=2

* INVx1_ASAP7_6t_L U26
MMN430_U26_inst39_MM0 y_4_ n42 VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MMP431_U26_inst39_MM1 y_4_ n42 VDD VDD pmos_lvt w=54.0n l=20n nfin=2

* INVx1_ASAP7_6t_L U27
MMN432_U27_inst40_MM0 n26 n41 VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MMP433_U27_inst40_MM1 n26 n41 VDD VDD pmos_lvt w=54.0n l=20n nfin=2

* INVx1_ASAP7_6t_L U28
MMN434_U28_inst41_MM0 y_3_ n40 VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MMP435_U28_inst41_MM1 y_3_ n40 VDD VDD pmos_lvt w=54.0n l=20n nfin=2

* INVx1_ASAP7_6t_L U29
MMN436_U29_inst42_MM0 n28 n39 VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MMP437_U29_inst42_MM1 n28 n39 VDD VDD pmos_lvt w=54.0n l=20n nfin=2

* INVx1_ASAP7_6t_L U30
MMN438_U30_inst43_MM0 y_2_ n38 VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MMP439_U30_inst43_MM1 y_2_ n38 VDD VDD pmos_lvt w=54.0n l=20n nfin=2

* INVx1_ASAP7_6t_L U31
MMN440_U31_inst44_MM0 n30 n37 VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MMP441_U31_inst44_MM1 n30 n37 VDD VDD pmos_lvt w=54.0n l=20n nfin=2

* INVx1_ASAP7_6t_L U32
MMN442_U32_inst45_MM0 y_1_ n36 VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MMP443_U32_inst45_MM1 y_1_ n36 VDD VDD pmos_lvt w=54.0n l=20n nfin=2

* INVx1_ASAP7_6t_L U33
MMN444_U33_inst46_MM0 n32 n35 VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MMP445_U33_inst46_MM1 n32 n35 VDD VDD pmos_lvt w=54.0n l=20n nfin=2

* INVx1_ASAP7_6t_L U34
MMN446_U34_inst47_MM0 y_0_ n34 VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MMP447_U34_inst47_MM1 y_0_ n34 VDD VDD pmos_lvt w=54.0n l=20n nfin=2

.ENDS
