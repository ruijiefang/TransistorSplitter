.SUBCKT ICGx1_ASAP7_75t_L CLK ENA GCLK SE VDD VSS
MM18 nos1 SE VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MM16 gclkn CLK VDD VDD pmos_lvt w=108.00n l=20n nfin=4
MM7 MS MH VDD VDD pmos_lvt w=27n l=20n nfin=1
MM11 pd2 MS VDD VDD pmos_lvt w=27n l=20n nfin=1
MM10 MH clkn pd2 VDD pmos_lvt w=27n l=20n nfin=1
MM1 MH CLK pu1 VDD pmos_lvt w=81.0n l=20n nfin=3
MM3 pu1 net0121 VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM21 clkn CLK VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM25 GCLK gclkn VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM26 net0121 ENA nos1 VDD pmos_lvt w=54.0n l=20n nfin=2
MM0 gclkn MH VDD VDD pmos_lvt w=108.00n l=20n nfin=4
MM2 gclkn CLK net0140 VSS nmos_lvt w=81.0n l=20n nfin=3
MM12 net0141 MH VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM14 net0140 MH VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM6 MS MH VSS VSS nmos_lvt w=27.0n l=20n nfin=1
MM13 gclkn CLK net0141 VSS nmos_lvt w=81.0n l=20n nfin=3
MM9 MH CLK pd3 VSS nmos_lvt w=27.0n l=20n nfin=1
MM8 pd3 MS VSS VSS nmos_lvt w=27.0n l=20n nfin=1
MM27 net0121 SE VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MM19 net0121 ENA VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MM24 GCLK gclkn VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM5 pd1 net0121 VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM4 MH clkn pd1 VSS nmos_lvt w=81.0n l=20n nfin=3
MM20 clkn CLK VSS VSS nmos_lvt w=81.0n l=20n nfin=3
.ENDS

