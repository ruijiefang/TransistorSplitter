.SUBCKT DFFLQNx1_ASAP7_75t_L CLK D QN VDD VSS
MM24 QN SH VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM23 clkb clkn VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MM20 clkn CLK VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MM17 SH clkb net0107 VSS nmos_lvt w=27.0n l=20n nfin=1
MM16 net0107 SS VSS VSS nmos_lvt w=27.0n l=20n nfin=1
MM14 SS SH VSS VSS nmos_lvt w=27.0n l=20n nfin=1
MM12 net029 clkn SH VSS nmos_lvt w=27.0n l=20n nfin=1
MM9 MH clkn net0109 VSS nmos_lvt w=27.0n l=20n nfin=1
MM8 net0109 net029 VSS VSS nmos_lvt w=27.0n l=20n nfin=1
MM6 net029 MH VSS VSS nmos_lvt w=27.0n l=20n nfin=1
MM5 net020 D VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM4 MH clkb net020 VSS nmos_lvt w=81.0n l=20n nfin=3
MM25 QN SH VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM13 net029 clkb SH VDD pmos_lvt w=27n l=20n nfin=1
MM22 clkb clkn VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MM21 clkn CLK VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MM19 net0108 SS VDD VDD pmos_lvt w=27.0n l=20n nfin=1
MM18 SH clkn net0108 VDD pmos_lvt w=27.0n l=20n nfin=1
MM15 SS SH VDD VDD pmos_lvt w=27.0n l=20n nfin=1
MM11 net0110 net029 VDD VDD pmos_lvt w=27.0n l=20n nfin=1
MM10 MH clkb net0110 VDD pmos_lvt w=27.0n l=20n nfin=1
MM7 net029 MH VDD VDD pmos_lvt w=27.0n l=20n nfin=1
MM1 MH clkn net06 VDD pmos_lvt w=81.0n l=20n nfin=3
MM3 net06 D VDD VDD pmos_lvt w=81.0n l=20n nfin=3
.ENDS

