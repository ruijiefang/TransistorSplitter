.SUBCKT ICGx2p67DC_ASAP7_75t_L CLK ENA GCLK SE VDD VSS
MM55 net0175 net0175 VDD VDD pmos_lvt w=162.00n l=20n nfin=6
MM54 net0175 net0212 VDD VDD pmos_lvt w=162.00n l=20n nfin=6
MM51 net0162 net0162 VDD VDD pmos_lvt w=162.00n l=20n nfin=6
MM47 gclkn2 CLK VDD VDD pmos_lvt w=108.00n l=20n nfin=4
MM46 gclkn2 MH VDD VDD pmos_lvt w=108.00n l=20n nfin=4
MM45 GCLK gclkn2 VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MM18 nos1 SE VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MM16 gclkn0 CLK VDD VDD pmos_lvt w=108.00n l=20n nfin=4
MM7 MS MH VDD VDD pmos_lvt w=27n l=20n nfin=1
MM11 pd2 MS VDD VDD pmos_lvt w=27n l=20n nfin=1
MM10 MH clkn pd2 VDD pmos_lvt w=27n l=20n nfin=1
MM25 GCLK gclkn0 VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MM50 net0162 net0207 VDD VDD pmos_lvt w=162.00n l=20n nfin=6
MM1 MH CLK pu1 VDD pmos_lvt w=81.0n l=20n nfin=3
MM3 pu1 net0121 VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM21 clkn CLK VDD VDD pmos_lvt w=162.00n l=20n nfin=6
MM29 GCLK gclkn1 VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MM30 gclkn1 MH VDD VDD pmos_lvt w=108.00n l=20n nfin=4
MM35 gclkn3 CLK VDD VDD pmos_lvt w=108.00n l=20n nfin=4
MM36 gclkn3 MH VDD VDD pmos_lvt w=108.00n l=20n nfin=4
MM37 GCLK gclkn3 VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MM31 gclkn1 CLK VDD VDD pmos_lvt w=108.00n l=20n nfin=4
MM26 net0121 ENA nos1 VDD pmos_lvt w=54.0n l=20n nfin=2
MM0 gclkn0 MH VDD VDD pmos_lvt w=108.00n l=20n nfin=4
MM57 net0212 net0175 VSS VSS nmos_lvt w=162.00n l=20n nfin=6
MM56 net0212 net0212 VSS VSS nmos_lvt w=162.00n l=20n nfin=6
MM53 net0207 net0162 VSS VSS nmos_lvt w=162.00n l=20n nfin=6
MM52 net0207 net0207 VSS VSS nmos_lvt w=162.00n l=20n nfin=6
MM27 net0121 SE VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MM13 gclkn0 CLK net0141 VSS nmos_lvt w=81.0n l=20n nfin=3
MM39 gclkn3 CLK net0244 VSS nmos_lvt w=81.0n l=20n nfin=3
MM6 MS MH VSS VSS nmos_lvt w=27.0n l=20n nfin=1
MM12 net0141 MH VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM40 net0243 MH VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM38 GCLK gclkn3 VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MM14 net0140 MH VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM2 gclkn0 CLK net0140 VSS nmos_lvt w=81.0n l=20n nfin=3
MM19 net0121 ENA VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MM9 MH CLK pd3 VSS nmos_lvt w=27.0n l=20n nfin=1
MM8 pd3 MS VSS VSS nmos_lvt w=27.0n l=20n nfin=1
MM15 net0247 MH VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM5 pd1 net0121 VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM4 MH clkn pd1 VSS nmos_lvt w=81.0n l=20n nfin=3
MM17 net0246 MH VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM22 gclkn1 CLK net0247 VSS nmos_lvt w=81.0n l=20n nfin=3
MM41 net0242 MH VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM42 gclkn2 CLK net0243 VSS nmos_lvt w=81.0n l=20n nfin=3
MM43 gclkn2 CLK net0242 VSS nmos_lvt w=81.0n l=20n nfin=3
MM32 net0245 MH VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM33 net0244 MH VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM20 clkn CLK VSS VSS nmos_lvt w=162.00n l=20n nfin=6
MM24 GCLK gclkn0 VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MM23 gclkn1 CLK net0246 VSS nmos_lvt w=81.0n l=20n nfin=3
MM34 gclkn3 CLK net0245 VSS nmos_lvt w=81.0n l=20n nfin=3
MM44 GCLK gclkn2 VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MM28 GCLK gclkn1 VSS VSS nmos_lvt w=54.0n l=20n nfin=2
.ENDS
