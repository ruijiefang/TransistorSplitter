.SUBCKT DLLx1_ASAP7_75t_L CLK D Q VDD VSS
MM23 clkb clkn VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MM5 pd1 D VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM4 MH clkn pd1 VSS nmos_lvt w=81.0n l=20n nfin=3
MM20 clkn CLK VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MM24 Q MH VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM6 net085 MH VSS VSS nmos_lvt w=27.0n l=20n nfin=1
MM9 MH clkb pd3 VSS nmos_lvt w=27.0n l=20n nfin=1
MM8 pd3 net085 VSS VSS nmos_lvt w=27.0n l=20n nfin=1
MM22 clkb clkn VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MM1 MH clkb pu1 VDD pmos_lvt w=81.0n l=20n nfin=3
MM3 pu1 D VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM25 Q MH VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM21 clkn CLK VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MM7 net085 MH VDD VDD pmos_lvt w=27n l=20n nfin=1
MM11 pd2 net085 VDD VDD pmos_lvt w=27n l=20n nfin=1
MM10 MH clkn pd2 VDD pmos_lvt w=27n l=20n nfin=1
.ENDS


.SUBCKT DLLx2_ASAP7_75t_L CLK D Q VDD VSS
MM23 clkb clkn VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MM5 pd1 D VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM4 MH clkn pd1 VSS nmos_lvt w=81.0n l=20n nfin=3
MM24 Q MH VSS VSS nmos_lvt w=162.00n l=20n nfin=6
MM20 clkn CLK VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MM6 net085 MH VSS VSS nmos_lvt w=27.0n l=20n nfin=1
MM9 MH clkb pd3 VSS nmos_lvt w=27.0n l=20n nfin=1
MM8 pd3 net085 VSS VSS nmos_lvt w=27.0n l=20n nfin=1
MM11 pd2 net085 VDD VDD pmos_lvt w=27n l=20n nfin=1
MM10 MH clkn pd2 VDD pmos_lvt w=27n l=20n nfin=1
MM22 clkb clkn VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MM1 MH clkb pu1 VDD pmos_lvt w=81.0n l=20n nfin=3
MM3 pu1 D VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM21 clkn CLK VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MM25 Q MH VDD VDD pmos_lvt w=162.00n l=20n nfin=6
MM7 net085 MH VDD VDD pmos_lvt w=27n l=20n nfin=1
.ENDS


.SUBCKT DLLx3_ASAP7_75t_L CLK D Q VDD VSS
MM24 Q MH VSS VSS nmos_lvt w=243.00n l=20n nfin=9
MM6 net30 MH VSS VSS nmos_lvt w=27.0n l=20n nfin=1
MM9 MH clkb pd3 VSS nmos_lvt w=27.0n l=20n nfin=1
MM8 pd3 net30 VSS VSS nmos_lvt w=27.0n l=20n nfin=1
MM23 clkb clkn VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MM5 pd1 D VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM4 MH clkn pd1 VSS nmos_lvt w=81.0n l=20n nfin=3
MM20 clkn CLK VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MM25 Q MH VDD VDD pmos_lvt w=243.00n l=20n nfin=9
MM7 net30 MH VDD VDD pmos_lvt w=27n l=20n nfin=1
MM11 pd2 net30 VDD VDD pmos_lvt w=27n l=20n nfin=1
MM10 MH clkn pd2 VDD pmos_lvt w=27n l=20n nfin=1
MM22 clkb clkn VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MM1 MH clkb pu1 VDD pmos_lvt w=81.0n l=20n nfin=3
MM3 pu1 D VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM21 clkn CLK VDD VDD pmos_lvt w=54.0n l=20n nfin=2
.ENDS


.SUBCKT FAx1_ASAP7_75t_L A B CI CON SN VDD VSS
MM22 SN CI net081 VDD pmos_lvt w=81.0n l=20n nfin=3
MM21 net081 B net082 VDD pmos_lvt w=81.0n l=20n nfin=3
MM20 net082 A VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM15 SN CON net027 VDD pmos_lvt w=81.0n l=20n nfin=3
MM14 net027 CI VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM13 net027 B VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM12 net027 A VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM5 CON A net37 VDD pmos_lvt w=81.0n l=20n nfin=3
MM6 net37 B VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM2 net27 B VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM1 CON CI net27 VDD pmos_lvt w=81.0n l=20n nfin=3
MM0 net27 A VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM25 SN CI net080 VSS nmos_lvt w=81.0n l=20n nfin=3
MM24 net080 B net079 VSS nmos_lvt w=81.0n l=20n nfin=3
MM23 net079 A VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM19 VSS CI net067 VSS nmos_lvt w=81.0n l=20n nfin=3
MM18 VSS B net067 VSS nmos_lvt w=81.0n l=20n nfin=3
MM17 VSS A net067 VSS nmos_lvt w=81.0n l=20n nfin=3
MM16 net067 CON SN VSS nmos_lvt w=81.0n l=20n nfin=3
MM11 VSS B net25 VSS nmos_lvt w=81.0n l=20n nfin=3
MM10 VSS B net36 VSS nmos_lvt w=81.0n l=20n nfin=3
MM9 VSS A net25 VSS nmos_lvt w=81.0n l=20n nfin=3
MM8 net36 A CON VSS nmos_lvt w=81.0n l=20n nfin=3
MM7 net25 CI CON VSS nmos_lvt w=81.0n l=20n nfin=3
.ENDS
